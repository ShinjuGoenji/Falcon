`ifdef RTL
    `define CYCLE_TIME 2.0
`endif
`ifdef GATE
    `define CYCLE_TIME 2.0
`endif

module PATTERN #(
    parameter   FLOAT_PRECISION = 64,
    parameter   logn = 8
)(
    // Output signals
    clk,
    rst_n,
    in_valid,
    fi_re, fi_im,
    s_re_1, s_im_1,
    s_re_2, s_im_2,
    s_re_3, s_im_3,
    s_re_4, s_im_4,
    s_re_5, s_im_5,
    s_re_6, s_im_6,
    s_re_7, s_im_7,
    s_re_8, s_im_8,
    // Input signals
    out_valid,
    tw_idx_1, 
    tw_idx_2, 
    tw_idx_3,
    tw_idx_4,
    tw_idx_5,
    tw_idx_6,
    tw_idx_7,
    tw_idx_8,
    fo_re, fo_im
);

parameter n = 1 << logn;

//---------------------------------------------------------------------
//   Input & Output
//---------------------------------------------------------------------
output reg                       clk;
output reg                       rst_n;
output reg                       in_valid;
output reg [FLOAT_PRECISION-1:0] fi_re;
output reg [FLOAT_PRECISION-1:0] fi_im;
output reg [FLOAT_PRECISION-1:0] s_re_1, s_im_1;
output reg [FLOAT_PRECISION-1:0] s_re_2, s_im_2;
output reg [FLOAT_PRECISION-1:0] s_re_3, s_im_3;
output reg [FLOAT_PRECISION-1:0] s_re_4, s_im_4;
output reg [FLOAT_PRECISION-1:0] s_re_5, s_im_5;
output reg [FLOAT_PRECISION-1:0] s_re_6, s_im_6;
output reg [FLOAT_PRECISION-1:0] s_re_7, s_im_7;
output reg [FLOAT_PRECISION-1:0] s_re_8, s_im_8;

input                  	 	out_valid;
input [logn:0]          	tw_idx_1;
input [logn:0]          	tw_idx_2;
input [logn:0]          	tw_idx_3;
input [logn:0]          	tw_idx_4;
input [logn:0]          	tw_idx_5;
input [logn:0]          	tw_idx_6;
input [logn:0]          	tw_idx_7;
input [logn:0]          	tw_idx_8;
input [FLOAT_PRECISION-1:0] fo_re;
input [FLOAT_PRECISION-1:0] fo_im;

//---------------------------------------------------------------------
//   Parameter & Integer
//---------------------------------------------------------------------
parameter INPUT_PATH  = "../00_TESTBED/input.txt";
parameter INDEX_PATH  = "../00_TESTBED/index.txt";
parameter OUTPUT_PATH = "../00_TESTBED/output8.txt";
parameter PATNUM_PATH = "../00_TESTBED/PATNUM.txt";
integer file_in, file_idx, file_out, file_num;

parameter MAX_OUT_LATENCY = 2000;
integer total_latency, out_latency, pattern_latency;
integer random_delay;

integer i_pat, i_in_deg, i_delay, i_out_deg;
integer PAT_NUM;

integer fscanf_int;

parameter [63:0] fpr_gm_tab [0:2047] = {
	64'h3ff0000000000000, 64'h0000000000000000,
	64'h8000000000000000, 64'h3ff0000000000000,
	64'h3fe6a09e667f3bcd, 64'h3fe6a09e667f3bcd,
	64'hbfe6a09e667f3bcd, 64'h3fe6a09e667f3bcd,
	64'h3fed906bcf328d46, 64'h3fd87de2a6aea963,
	64'hbfd87de2a6aea963, 64'h3fed906bcf328d46,
	64'h3fd87de2a6aea963, 64'h3fed906bcf328d46,
	64'hbfed906bcf328d46, 64'h3fd87de2a6aea963,
	64'h3fef6297cff75cb0, 64'h3fc8f8b83c69a60b,
	64'hbfc8f8b83c69a60b, 64'h3fef6297cff75cb0,
	64'h3fe1c73b39ae68c8, 64'h3fea9b66290ea1a3,
	64'hbfea9b66290ea1a3, 64'h3fe1c73b39ae68c8,
	64'h3fea9b66290ea1a3, 64'h3fe1c73b39ae68c8,
	64'hbfe1c73b39ae68c8, 64'h3fea9b66290ea1a3,
	64'h3fc8f8b83c69a60b, 64'h3fef6297cff75cb0,
	64'hbfef6297cff75cb0, 64'h3fc8f8b83c69a60b,
	64'h3fefd88da3d12526, 64'h3fb917a6bc29b42c,
	64'hbfb917a6bc29b42c, 64'h3fefd88da3d12526,
	64'h3fe44cf325091dd6, 64'h3fe8bc806b151741,
	64'hbfe8bc806b151741, 64'h3fe44cf325091dd6,
	64'h3fec38b2f180bdb1, 64'h3fde2b5d3806f63b,
	64'hbfde2b5d3806f63b, 64'h3fec38b2f180bdb1,
	64'h3fd294062ed59f06, 64'h3fee9f4156c62dda,
	64'hbfee9f4156c62dda, 64'h3fd294062ed59f06,
	64'h3fee9f4156c62dda, 64'h3fd294062ed59f06,
	64'hbfd294062ed59f06, 64'h3fee9f4156c62dda,
	64'h3fde2b5d3806f63b, 64'h3fec38b2f180bdb1,
	64'hbfec38b2f180bdb1, 64'h3fde2b5d3806f63b,
	64'h3fe8bc806b151741, 64'h3fe44cf325091dd6,
	64'hbfe44cf325091dd6, 64'h3fe8bc806b151741,
	64'h3fb917a6bc29b42c, 64'h3fefd88da3d12526,
	64'hbfefd88da3d12526, 64'h3fb917a6bc29b42c,
	64'h3feff621e3796d7e, 64'h3fa91f65f10dd814,
	64'hbfa91f65f10dd814, 64'h3feff621e3796d7e,
	64'h3fe57d69348ceca0, 64'h3fe7b5df226aafaf,
	64'hbfe7b5df226aafaf, 64'h3fe57d69348ceca0,
	64'h3feced7af43cc773, 64'h3fdb5d1009e15cc0,
	64'hbfdb5d1009e15cc0, 64'h3feced7af43cc773,
	64'h3fd58f9a75ab1fdd, 64'h3fee212104f686e5,
	64'hbfee212104f686e5, 64'h3fd58f9a75ab1fdd,
	64'h3fef0a7efb9230d7, 64'h3fcf19f97b215f1b,
	64'hbfcf19f97b215f1b, 64'h3fef0a7efb9230d7,
	64'h3fe073879922ffee, 64'h3feb728345196e3e,
	64'hbfeb728345196e3e, 64'h3fe073879922ffee,
	64'h3fe9b3e047f38741, 64'h3fe30ff7fce17035,
	64'hbfe30ff7fce17035, 64'h3fe9b3e047f38741,
	64'h3fc2c8106e8e613a, 64'h3fefa7557f08a517,
	64'hbfefa7557f08a517, 64'h3fc2c8106e8e613a,
	64'h3fefa7557f08a517, 64'h3fc2c8106e8e613a,
	64'hbfc2c8106e8e613a, 64'h3fefa7557f08a517,
	64'h3fe30ff7fce17035, 64'h3fe9b3e047f38741,
	64'hbfe9b3e047f38741, 64'h3fe30ff7fce17035,
	64'h3feb728345196e3e, 64'h3fe073879922ffee,
	64'hbfe073879922ffee, 64'h3feb728345196e3e,
	64'h3fcf19f97b215f1b, 64'h3fef0a7efb9230d7,
	64'hbfef0a7efb9230d7, 64'h3fcf19f97b215f1b,
	64'h3fee212104f686e5, 64'h3fd58f9a75ab1fdd,
	64'hbfd58f9a75ab1fdd, 64'h3fee212104f686e5,
	64'h3fdb5d1009e15cc0, 64'h3feced7af43cc773,
	64'hbfeced7af43cc773, 64'h3fdb5d1009e15cc0,
	64'h3fe7b5df226aafaf, 64'h3fe57d69348ceca0,
	64'hbfe57d69348ceca0, 64'h3fe7b5df226aafaf,
	64'h3fa91f65f10dd814, 64'h3feff621e3796d7e,
	64'hbfeff621e3796d7e, 64'h3fa91f65f10dd814,
	64'h3feffd886084cd0d, 64'h3f992155f7a3667e,
	64'hbf992155f7a3667e, 64'h3feffd886084cd0d,
	64'h3fe610b7551d2cdf, 64'h3fe72d0837efff96,
	64'hbfe72d0837efff96, 64'h3fe610b7551d2cdf,
	64'h3fed4134d14dc93a, 64'h3fd9ef7943a8ed8a,
	64'hbfd9ef7943a8ed8a, 64'h3fed4134d14dc93a,
	64'h3fd7088530fa459f, 64'h3feddb13b6ccc23c,
	64'hbfeddb13b6ccc23c, 64'h3fd7088530fa459f,
	64'h3fef38f3ac64e589, 64'h3fcc0b826a7e4f63,
	64'hbfcc0b826a7e4f63, 64'h3fef38f3ac64e589,
	64'h3fe11eb3541b4b23, 64'h3feb090a58150200,
	64'hbfeb090a58150200, 64'h3fe11eb3541b4b23,
	64'h3fea29a7a0462782, 64'h3fe26d054cdd12df,
	64'hbfe26d054cdd12df, 64'h3fea29a7a0462782,
	64'h3fc5e214448b3fc6, 64'h3fef8764fa714ba9,
	64'hbfef8764fa714ba9, 64'h3fc5e214448b3fc6,
	64'h3fefc26470e19fd3, 64'h3fbf564e56a9730e,
	64'hbfbf564e56a9730e, 64'h3fefc26470e19fd3,
	64'h3fe3affa292050b9, 64'h3fe93a22499263fb,
	64'hbfe93a22499263fb, 64'h3fe3affa292050b9,
	64'h3febd7c0ac6f952a, 64'h3fdf8ba4dbf89aba,
	64'hbfdf8ba4dbf89aba, 64'h3febd7c0ac6f952a,
	64'h3fd111d262b1f677, 64'h3feed740e7684963,
	64'hbfeed740e7684963, 64'h3fd111d262b1f677,
	64'h3fee6288ec48e112, 64'h3fd4135c94176601,
	64'hbfd4135c94176601, 64'h3fee6288ec48e112,
	64'h3fdcc66e9931c45e, 64'h3fec954b213411f5,
	64'hbfec954b213411f5, 64'h3fdcc66e9931c45e,
	64'h3fe83b0e0bff976e, 64'h3fe4e6cabbe3e5e9,
	64'hbfe4e6cabbe3e5e9, 64'h3fe83b0e0bff976e,
	64'h3fb2d52092ce19f6, 64'h3fefe9cdad01883a,
	64'hbfefe9cdad01883a, 64'h3fb2d52092ce19f6,
	64'h3fefe9cdad01883a, 64'h3fb2d52092ce19f6,
	64'hbfb2d52092ce19f6, 64'h3fefe9cdad01883a,
	64'h3fe4e6cabbe3e5e9, 64'h3fe83b0e0bff976e,
	64'hbfe83b0e0bff976e, 64'h3fe4e6cabbe3e5e9,
	64'h3fec954b213411f5, 64'h3fdcc66e9931c45e,
	64'hbfdcc66e9931c45e, 64'h3fec954b213411f5,
	64'h3fd4135c94176601, 64'h3fee6288ec48e112,
	64'hbfee6288ec48e112, 64'h3fd4135c94176601,
	64'h3feed740e7684963, 64'h3fd111d262b1f677,
	64'hbfd111d262b1f677, 64'h3feed740e7684963,
	64'h3fdf8ba4dbf89aba, 64'h3febd7c0ac6f952a,
	64'hbfebd7c0ac6f952a, 64'h3fdf8ba4dbf89aba,
	64'h3fe93a22499263fb, 64'h3fe3affa292050b9,
	64'hbfe3affa292050b9, 64'h3fe93a22499263fb,
	64'h3fbf564e56a9730e, 64'h3fefc26470e19fd3,
	64'hbfefc26470e19fd3, 64'h3fbf564e56a9730e,
	64'h3fef8764fa714ba9, 64'h3fc5e214448b3fc6,
	64'hbfc5e214448b3fc6, 64'h3fef8764fa714ba9,
	64'h3fe26d054cdd12df, 64'h3fea29a7a0462782,
	64'hbfea29a7a0462782, 64'h3fe26d054cdd12df,
	64'h3feb090a58150200, 64'h3fe11eb3541b4b23,
	64'hbfe11eb3541b4b23, 64'h3feb090a58150200,
	64'h3fcc0b826a7e4f63, 64'h3fef38f3ac64e589,
	64'hbfef38f3ac64e589, 64'h3fcc0b826a7e4f63,
	64'h3feddb13b6ccc23c, 64'h3fd7088530fa459f,
	64'hbfd7088530fa459f, 64'h3feddb13b6ccc23c,
	64'h3fd9ef7943a8ed8a, 64'h3fed4134d14dc93a,
	64'hbfed4134d14dc93a, 64'h3fd9ef7943a8ed8a,
	64'h3fe72d0837efff96, 64'h3fe610b7551d2cdf,
	64'hbfe610b7551d2cdf, 64'h3fe72d0837efff96,
	64'h3f992155f7a3667e, 64'h3feffd886084cd0d,
	64'hbfeffd886084cd0d, 64'h3f992155f7a3667e,
	64'h3fefff62169b92db, 64'h3f8921d1fcdec784,
	64'hbf8921d1fcdec784, 64'h3fefff62169b92db,
	64'h3fe6591925f0783d, 64'h3fe6e74454eaa8af,
	64'hbfe6e74454eaa8af, 64'h3fe6591925f0783d,
	64'h3fed696173c9e68b, 64'h3fd9372a63bc93d7,
	64'hbfd9372a63bc93d7, 64'h3fed696173c9e68b,
	64'h3fd7c3a9311dcce7, 64'h3fedb6526238a09b,
	64'hbfedb6526238a09b, 64'h3fd7c3a9311dcce7,
	64'h3fef4e603b0b2f2d, 64'h3fca82a025b00451,
	64'hbfca82a025b00451, 64'h3fef4e603b0b2f2d,
	64'h3fe1734d63dedb49, 64'h3fead2bc9e21d511,
	64'hbfead2bc9e21d511, 64'h3fe1734d63dedb49,
	64'h3fea63091b02fae2, 64'h3fe21a799933eb59,
	64'hbfe21a799933eb59, 64'h3fea63091b02fae2,
	64'h3fc76dd9de50bf31, 64'h3fef7599a3a12077,
	64'hbfef7599a3a12077, 64'h3fc76dd9de50bf31,
	64'h3fefce15fd6da67b, 64'h3fbc3785c79ec2d5,
	64'hbfbc3785c79ec2d5, 64'h3fefce15fd6da67b,
	64'h3fe3fed9534556d4, 64'h3fe8fbcca3ef940d,
	64'hbfe8fbcca3ef940d, 64'h3fe3fed9534556d4,
	64'h3fec08c426725549, 64'h3fdedc1952ef78d6,
	64'hbfdedc1952ef78d6, 64'h3fec08c426725549,
	64'h3fd1d3443f4cdb3e, 64'h3feebbd8c8df0b74,
	64'hbfeebbd8c8df0b74, 64'h3fd1d3443f4cdb3e,
	64'h3fee817bab4cd10d, 64'h3fd35410c2e18152,
	64'hbfd35410c2e18152, 64'h3fee817bab4cd10d,
	64'h3fdd79775b86e389, 64'h3fec678b3488739b,
	64'hbfec678b3488739b, 64'h3fdd79775b86e389,
	64'h3fe87c400fba2ebf, 64'h3fe49a449b9b0939,
	64'hbfe49a449b9b0939, 64'h3fe87c400fba2ebf,
	64'h3fb5f6d00a9aa419, 64'h3fefe1cafcbd5b09,
	64'hbfefe1cafcbd5b09, 64'h3fb5f6d00a9aa419,
	64'h3feff095658e71ad, 64'h3faf656e79f820e0,
	64'hbfaf656e79f820e0, 64'h3feff095658e71ad,
	64'h3fe5328292a35596, 64'h3fe7f8ece3571771,
	64'hbfe7f8ece3571771, 64'h3fe5328292a35596,
	64'h3fecc1f0f3fcfc5c, 64'h3fdc1249d8011ee7,
	64'hbfdc1249d8011ee7, 64'h3fecc1f0f3fcfc5c,
	64'h3fd4d1e24278e76a, 64'h3fee426a4b2bc17e,
	64'hbfee426a4b2bc17e, 64'h3fd4d1e24278e76a,
	64'h3feef178a3e473c2, 64'h3fd04fb80e37fdae,
	64'hbfd04fb80e37fdae, 64'h3feef178a3e473c2,
	64'h3fe01cfc874c3eb7, 64'h3feba5aa673590d2,
	64'hbfeba5aa673590d2, 64'h3fe01cfc874c3eb7,
	64'h3fe9777ef4c7d742, 64'h3fe36058b10659f3,
	64'hbfe36058b10659f3, 64'h3fe9777ef4c7d742,
	64'h3fc139f0cedaf577, 64'h3fefb5797195d741,
	64'hbfefb5797195d741, 64'h3fc139f0cedaf577,
	64'h3fef97f924c9099b, 64'h3fc45576b1293e5a,
	64'hbfc45576b1293e5a, 64'h3fef97f924c9099b,
	64'h3fe2bedb25faf3ea, 64'h3fe9ef43ef29af94,
	64'hbfe9ef43ef29af94, 64'h3fe2bedb25faf3ea,
	64'h3feb3e4d3ef55712, 64'h3fe0c9704d5d898f,
	64'hbfe0c9704d5d898f, 64'h3feb3e4d3ef55712,
	64'h3fcd934fe5454311, 64'h3fef2252f7763ada,
	64'hbfef2252f7763ada, 64'h3fcd934fe5454311,
	64'h3fedfeae622dbe2b, 64'h3fd64c7ddd3f27c6,
	64'hbfd64c7ddd3f27c6, 64'h3fedfeae622dbe2b,
	64'h3fdaa6c82b6d3fca, 64'h3fed17e7743e35dc,
	64'hbfed17e7743e35dc, 64'h3fdaa6c82b6d3fca,
	64'h3fe771e75f037261, 64'h3fe5c77bbe65018c,
	64'hbfe5c77bbe65018c, 64'h3fe771e75f037261,
	64'h3fa2d865759455cd, 64'h3feffa72effef75d,
	64'hbfeffa72effef75d, 64'h3fa2d865759455cd,
	64'h3feffa72effef75d, 64'h3fa2d865759455cd,
	64'hbfa2d865759455cd, 64'h3feffa72effef75d,
	64'h3fe5c77bbe65018c, 64'h3fe771e75f037261,
	64'hbfe771e75f037261, 64'h3fe5c77bbe65018c,
	64'h3fed17e7743e35dc, 64'h3fdaa6c82b6d3fca,
	64'hbfdaa6c82b6d3fca, 64'h3fed17e7743e35dc,
	64'h3fd64c7ddd3f27c6, 64'h3fedfeae622dbe2b,
	64'hbfedfeae622dbe2b, 64'h3fd64c7ddd3f27c6,
	64'h3fef2252f7763ada, 64'h3fcd934fe5454311,
	64'hbfcd934fe5454311, 64'h3fef2252f7763ada,
	64'h3fe0c9704d5d898f, 64'h3feb3e4d3ef55712,
	64'hbfeb3e4d3ef55712, 64'h3fe0c9704d5d898f,
	64'h3fe9ef43ef29af94, 64'h3fe2bedb25faf3ea,
	64'hbfe2bedb25faf3ea, 64'h3fe9ef43ef29af94,
	64'h3fc45576b1293e5a, 64'h3fef97f924c9099b,
	64'hbfef97f924c9099b, 64'h3fc45576b1293e5a,
	64'h3fefb5797195d741, 64'h3fc139f0cedaf577,
	64'hbfc139f0cedaf577, 64'h3fefb5797195d741,
	64'h3fe36058b10659f3, 64'h3fe9777ef4c7d742,
	64'hbfe9777ef4c7d742, 64'h3fe36058b10659f3,
	64'h3feba5aa673590d2, 64'h3fe01cfc874c3eb7,
	64'hbfe01cfc874c3eb7, 64'h3feba5aa673590d2,
	64'h3fd04fb80e37fdae, 64'h3feef178a3e473c2,
	64'hbfeef178a3e473c2, 64'h3fd04fb80e37fdae,
	64'h3fee426a4b2bc17e, 64'h3fd4d1e24278e76a,
	64'hbfd4d1e24278e76a, 64'h3fee426a4b2bc17e,
	64'h3fdc1249d8011ee7, 64'h3fecc1f0f3fcfc5c,
	64'hbfecc1f0f3fcfc5c, 64'h3fdc1249d8011ee7,
	64'h3fe7f8ece3571771, 64'h3fe5328292a35596,
	64'hbfe5328292a35596, 64'h3fe7f8ece3571771,
	64'h3faf656e79f820e0, 64'h3feff095658e71ad,
	64'hbfeff095658e71ad, 64'h3faf656e79f820e0,
	64'h3fefe1cafcbd5b09, 64'h3fb5f6d00a9aa419,
	64'hbfb5f6d00a9aa419, 64'h3fefe1cafcbd5b09,
	64'h3fe49a449b9b0939, 64'h3fe87c400fba2ebf,
	64'hbfe87c400fba2ebf, 64'h3fe49a449b9b0939,
	64'h3fec678b3488739b, 64'h3fdd79775b86e389,
	64'hbfdd79775b86e389, 64'h3fec678b3488739b,
	64'h3fd35410c2e18152, 64'h3fee817bab4cd10d,
	64'hbfee817bab4cd10d, 64'h3fd35410c2e18152,
	64'h3feebbd8c8df0b74, 64'h3fd1d3443f4cdb3e,
	64'hbfd1d3443f4cdb3e, 64'h3feebbd8c8df0b74,
	64'h3fdedc1952ef78d6, 64'h3fec08c426725549,
	64'hbfec08c426725549, 64'h3fdedc1952ef78d6,
	64'h3fe8fbcca3ef940d, 64'h3fe3fed9534556d4,
	64'hbfe3fed9534556d4, 64'h3fe8fbcca3ef940d,
	64'h3fbc3785c79ec2d5, 64'h3fefce15fd6da67b,
	64'hbfefce15fd6da67b, 64'h3fbc3785c79ec2d5,
	64'h3fef7599a3a12077, 64'h3fc76dd9de50bf31,
	64'hbfc76dd9de50bf31, 64'h3fef7599a3a12077,
	64'h3fe21a799933eb59, 64'h3fea63091b02fae2,
	64'hbfea63091b02fae2, 64'h3fe21a799933eb59,
	64'h3fead2bc9e21d511, 64'h3fe1734d63dedb49,
	64'hbfe1734d63dedb49, 64'h3fead2bc9e21d511,
	64'h3fca82a025b00451, 64'h3fef4e603b0b2f2d,
	64'hbfef4e603b0b2f2d, 64'h3fca82a025b00451,
	64'h3fedb6526238a09b, 64'h3fd7c3a9311dcce7,
	64'hbfd7c3a9311dcce7, 64'h3fedb6526238a09b,
	64'h3fd9372a63bc93d7, 64'h3fed696173c9e68b,
	64'hbfed696173c9e68b, 64'h3fd9372a63bc93d7,
	64'h3fe6e74454eaa8af, 64'h3fe6591925f0783d,
	64'hbfe6591925f0783d, 64'h3fe6e74454eaa8af,
	64'h3f8921d1fcdec784, 64'h3fefff62169b92db,
	64'hbfefff62169b92db, 64'h3f8921d1fcdec784,
	64'h3fefffd8858e8a92, 64'h3f7921f0fe670071,
	64'hbf7921f0fe670071, 64'h3fefffd8858e8a92,
	64'h3fe67cf78491af10, 64'h3fe6c40d73c18275,
	64'hbfe6c40d73c18275, 64'h3fe67cf78491af10,
	64'h3fed7d0b02b8ecf9, 64'h3fd8daa52ec8a4b0,
	64'hbfd8daa52ec8a4b0, 64'h3fed7d0b02b8ecf9,
	64'h3fd820e3b04eaac4, 64'h3feda383a9668988,
	64'hbfeda383a9668988, 64'h3fd820e3b04eaac4,
	64'h3fef58a2b1789e84, 64'h3fc9bdcbf2dc4366,
	64'hbfc9bdcbf2dc4366, 64'h3fef58a2b1789e84,
	64'h3fe19d5a09f2b9b8, 64'h3feab7325916c0d4,
	64'hbfeab7325916c0d4, 64'h3fe19d5a09f2b9b8,
	64'h3fea7f58529fe69d, 64'h3fe1f0f08bbc861b,
	64'hbfe1f0f08bbc861b, 64'h3fea7f58529fe69d,
	64'h3fc83366e89c64c6, 64'h3fef6c3f7df5bbb7,
	64'hbfef6c3f7df5bbb7, 64'h3fc83366e89c64c6,
	64'h3fefd37914220b84, 64'h3fbaa7b724495c03,
	64'hbfbaa7b724495c03, 64'h3fefd37914220b84,
	64'h3fe425ff178e6bb1, 64'h3fe8dc45331698cc,
	64'hbfe8dc45331698cc, 64'h3fe425ff178e6bb1,
	64'h3fec20de3fa971b0, 64'h3fde83e0eaf85114,
	64'hbfde83e0eaf85114, 64'h3fec20de3fa971b0,
	64'h3fd233bbabc3bb71, 64'h3feeadb2e8e7a88e,
	64'hbfeeadb2e8e7a88e, 64'h3fd233bbabc3bb71,
	64'h3fee9084361df7f2, 64'h3fd2f422daec0387,
	64'hbfd2f422daec0387, 64'h3fee9084361df7f2,
	64'h3fddd28f1481cc58, 64'h3fec5042012b6907,
	64'hbfec5042012b6907, 64'h3fddd28f1481cc58,
	64'h3fe89c7e9a4dd4aa, 64'h3fe473b51b987347,
	64'hbfe473b51b987347, 64'h3fe89c7e9a4dd4aa,
	64'h3fb787586a5d5b21, 64'h3fefdd539ff1f456,
	64'hbfefdd539ff1f456, 64'h3fb787586a5d5b21,
	64'h3feff3830f8d575c, 64'h3fac428d12c0d7e3,
	64'hbfac428d12c0d7e3, 64'h3feff3830f8d575c,
	64'h3fe5581038975137, 64'h3fe7d7836cc33db2,
	64'hbfe7d7836cc33db2, 64'h3fe5581038975137,
	64'h3fecd7d9898b32f6, 64'h3fdbb7cf2304bd01,
	64'hbfdbb7cf2304bd01, 64'h3fecd7d9898b32f6,
	64'h3fd530d880af3c24, 64'h3fee31eae870ce25,
	64'hbfee31eae870ce25, 64'h3fd530d880af3c24,
	64'h3feefe220c0b95ec, 64'h3fcfdcdc1adfedf9,
	64'hbfcfdcdc1adfedf9, 64'h3feefe220c0b95ec,
	64'h3fe0485626ae221a, 64'h3feb8c38d27504e9,
	64'hbfeb8c38d27504e9, 64'h3fe0485626ae221a,
	64'h3fe995cf2ed80d22, 64'h3fe338400d0c8e57,
	64'hbfe338400d0c8e57, 64'h3fe995cf2ed80d22,
	64'h3fc20116d4ec7bcf, 64'h3fefae8e8e46cfbb,
	64'hbfefae8e8e46cfbb, 64'h3fc20116d4ec7bcf,
	64'h3fef9fce55adb2c8, 64'h3fc38edbb0cd8d14,
	64'hbfc38edbb0cd8d14, 64'h3fef9fce55adb2c8,
	64'h3fe2e780e3e8ea17, 64'h3fe9d1b1f5ea80d5,
	64'hbfe9d1b1f5ea80d5, 64'h3fe2e780e3e8ea17,
	64'h3feb5889fe921405, 64'h3fe09e907417c5e1,
	64'hbfe09e907417c5e1, 64'h3feb5889fe921405,
	64'h3fce56ca1e101a1b, 64'h3fef168f53f7205d,
	64'hbfef168f53f7205d, 64'h3fce56ca1e101a1b,
	64'h3fee100cca2980ac, 64'h3fd5ee27379ea693,
	64'hbfd5ee27379ea693, 64'h3fee100cca2980ac,
	64'h3fdb020d6c7f4009, 64'h3fed02d4feb2bd92,
	64'hbfed02d4feb2bd92, 64'h3fdb020d6c7f4009,
	64'h3fe79400574f55e5, 64'h3fe5a28d2a5d7250,
	64'hbfe5a28d2a5d7250, 64'h3fe79400574f55e5,
	64'h3fa5fc00d290cd43, 64'h3feff871dadb81df,
	64'hbfeff871dadb81df, 64'h3fa5fc00d290cd43,
	64'h3feffc251df1d3f8, 64'h3f9f693731d1cf01,
	64'hbf9f693731d1cf01, 64'h3feffc251df1d3f8,
	64'h3fe5ec3495837074, 64'h3fe74f948da8d28d,
	64'hbfe74f948da8d28d, 64'h3fe5ec3495837074,
	64'h3fed2cb220e0ef9f, 64'h3fda4b4127dea1e5,
	64'hbfda4b4127dea1e5, 64'h3fed2cb220e0ef9f,
	64'h3fd6aa9d7dc77e17, 64'h3feded05f7de47da,
	64'hbfeded05f7de47da, 64'h3fd6aa9d7dc77e17,
	64'h3fef2dc9c9089a9d, 64'h3fcccf8cb312b286,
	64'hbfcccf8cb312b286, 64'h3fef2dc9c9089a9d,
	64'h3fe0f426bb2a8e7e, 64'h3feb23cd470013b4,
	64'hbfeb23cd470013b4, 64'h3fe0f426bb2a8e7e,
	64'h3fea0c95eabaf937, 64'h3fe2960727629ca8,
	64'hbfe2960727629ca8, 64'h3fea0c95eabaf937,
	64'h3fc51bdf8597c5f2, 64'h3fef8fd5ffae41db,
	64'hbfef8fd5ffae41db, 64'h3fc51bdf8597c5f2,
	64'h3fefbc1617e44186, 64'h3fc072a047ba831d,
	64'hbfc072a047ba831d, 64'h3fefbc1617e44186,
	64'h3fe3884185dfeb22, 64'h3fe958efe48e6dd7,
	64'hbfe958efe48e6dd7, 64'h3fe3884185dfeb22,
	64'h3febbed7c49380ea, 64'h3fdfe2f64be71210,
	64'hbfdfe2f64be71210, 64'h3febbed7c49380ea,
	64'h3fd0b0d9cfdbdb90, 64'h3feee482e25a9dbc,
	64'hbfeee482e25a9dbc, 64'h3fd0b0d9cfdbdb90,
	64'h3fee529f04729ffc, 64'h3fd472b8a5571054,
	64'hbfd472b8a5571054, 64'h3fee529f04729ffc,
	64'h3fdc6c7f4997000b, 64'h3fecabc169a0b900,
	64'hbfecabc169a0b900, 64'h3fdc6c7f4997000b,
	64'h3fe81a1b33b57acc, 64'h3fe50cc09f59a09b,
	64'hbfe50cc09f59a09b, 64'h3fe81a1b33b57acc,
	64'h3fb1440134d709b3, 64'h3fefed58ecb673c4,
	64'hbfefed58ecb673c4, 64'h3fb1440134d709b3,
	64'h3fefe5f3af2e3940, 64'h3fb4661179272096,
	64'hbfb4661179272096, 64'h3fefe5f3af2e3940,
	64'h3fe4c0a145ec0004, 64'h3fe85bc51ae958cc,
	64'hbfe85bc51ae958cc, 64'h3fe4c0a145ec0004,
	64'h3fec7e8e52233cf3, 64'h3fdd2016e8e9db5b,
	64'hbfdd2016e8e9db5b, 64'h3fec7e8e52233cf3,
	64'h3fd3b3cefa0414b7, 64'h3fee7227db6a9744,
	64'hbfee7227db6a9744, 64'h3fd3b3cefa0414b7,
	64'h3feec9b2d3c3bf84, 64'h3fd172a0d7765177,
	64'hbfd172a0d7765177, 64'h3feec9b2d3c3bf84,
	64'h3fdf3405963fd067, 64'h3febf064e15377dd,
	64'hbfebf064e15377dd, 64'h3fdf3405963fd067,
	64'h3fe91b166fd49da2, 64'h3fe3d78238c58344,
	64'hbfe3d78238c58344, 64'h3fe91b166fd49da2,
	64'h3fbdc70ecbae9fc9, 64'h3fefc8646cfeb721,
	64'hbfefc8646cfeb721, 64'h3fbdc70ecbae9fc9,
	64'h3fef7ea629e63d6e, 64'h3fc6a81304f64ab2,
	64'hbfc6a81304f64ab2, 64'h3fef7ea629e63d6e,
	64'h3fe243d5fb98ac1f, 64'h3fea4678c8119ac8,
	64'hbfea4678c8119ac8, 64'h3fe243d5fb98ac1f,
	64'h3feaee04b43c1474, 64'h3fe14915af336ceb,
	64'hbfe14915af336ceb, 64'h3feaee04b43c1474,
	64'h3fcb4732ef3d6722, 64'h3fef43d085ff92dd,
	64'hbfef43d085ff92dd, 64'h3fcb4732ef3d6722,
	64'h3fedc8d7cb410260, 64'h3fd766340f2418f6,
	64'hbfd766340f2418f6, 64'h3fedc8d7cb410260,
	64'h3fd993716141bdff, 64'h3fed556f52e93eb1,
	64'hbfed556f52e93eb1, 64'h3fd993716141bdff,
	64'h3fe70a42b3176d7a, 64'h3fe63503a31c1be9,
	64'hbfe63503a31c1be9, 64'h3fe70a42b3176d7a,
	64'h3f92d936bbe30efd, 64'h3feffe9cb44b51a1,
	64'hbfeffe9cb44b51a1, 64'h3f92d936bbe30efd,
	64'h3feffe9cb44b51a1, 64'h3f92d936bbe30efd,
	64'hbf92d936bbe30efd, 64'h3feffe9cb44b51a1,
	64'h3fe63503a31c1be9, 64'h3fe70a42b3176d7a,
	64'hbfe70a42b3176d7a, 64'h3fe63503a31c1be9,
	64'h3fed556f52e93eb1, 64'h3fd993716141bdff,
	64'hbfd993716141bdff, 64'h3fed556f52e93eb1,
	64'h3fd766340f2418f6, 64'h3fedc8d7cb410260,
	64'hbfedc8d7cb410260, 64'h3fd766340f2418f6,
	64'h3fef43d085ff92dd, 64'h3fcb4732ef3d6722,
	64'hbfcb4732ef3d6722, 64'h3fef43d085ff92dd,
	64'h3fe14915af336ceb, 64'h3feaee04b43c1474,
	64'hbfeaee04b43c1474, 64'h3fe14915af336ceb,
	64'h3fea4678c8119ac8, 64'h3fe243d5fb98ac1f,
	64'hbfe243d5fb98ac1f, 64'h3fea4678c8119ac8,
	64'h3fc6a81304f64ab2, 64'h3fef7ea629e63d6e,
	64'hbfef7ea629e63d6e, 64'h3fc6a81304f64ab2,
	64'h3fefc8646cfeb721, 64'h3fbdc70ecbae9fc9,
	64'hbfbdc70ecbae9fc9, 64'h3fefc8646cfeb721,
	64'h3fe3d78238c58344, 64'h3fe91b166fd49da2,
	64'hbfe91b166fd49da2, 64'h3fe3d78238c58344,
	64'h3febf064e15377dd, 64'h3fdf3405963fd067,
	64'hbfdf3405963fd067, 64'h3febf064e15377dd,
	64'h3fd172a0d7765177, 64'h3feec9b2d3c3bf84,
	64'hbfeec9b2d3c3bf84, 64'h3fd172a0d7765177,
	64'h3fee7227db6a9744, 64'h3fd3b3cefa0414b7,
	64'hbfd3b3cefa0414b7, 64'h3fee7227db6a9744,
	64'h3fdd2016e8e9db5b, 64'h3fec7e8e52233cf3,
	64'hbfec7e8e52233cf3, 64'h3fdd2016e8e9db5b,
	64'h3fe85bc51ae958cc, 64'h3fe4c0a145ec0004,
	64'hbfe4c0a145ec0004, 64'h3fe85bc51ae958cc,
	64'h3fb4661179272096, 64'h3fefe5f3af2e3940,
	64'hbfefe5f3af2e3940, 64'h3fb4661179272096,
	64'h3fefed58ecb673c4, 64'h3fb1440134d709b3,
	64'hbfb1440134d709b3, 64'h3fefed58ecb673c4,
	64'h3fe50cc09f59a09b, 64'h3fe81a1b33b57acc,
	64'hbfe81a1b33b57acc, 64'h3fe50cc09f59a09b,
	64'h3fecabc169a0b900, 64'h3fdc6c7f4997000b,
	64'hbfdc6c7f4997000b, 64'h3fecabc169a0b900,
	64'h3fd472b8a5571054, 64'h3fee529f04729ffc,
	64'hbfee529f04729ffc, 64'h3fd472b8a5571054,
	64'h3feee482e25a9dbc, 64'h3fd0b0d9cfdbdb90,
	64'hbfd0b0d9cfdbdb90, 64'h3feee482e25a9dbc,
	64'h3fdfe2f64be71210, 64'h3febbed7c49380ea,
	64'hbfebbed7c49380ea, 64'h3fdfe2f64be71210,
	64'h3fe958efe48e6dd7, 64'h3fe3884185dfeb22,
	64'hbfe3884185dfeb22, 64'h3fe958efe48e6dd7,
	64'h3fc072a047ba831d, 64'h3fefbc1617e44186,
	64'hbfefbc1617e44186, 64'h3fc072a047ba831d,
	64'h3fef8fd5ffae41db, 64'h3fc51bdf8597c5f2,
	64'hbfc51bdf8597c5f2, 64'h3fef8fd5ffae41db,
	64'h3fe2960727629ca8, 64'h3fea0c95eabaf937,
	64'hbfea0c95eabaf937, 64'h3fe2960727629ca8,
	64'h3feb23cd470013b4, 64'h3fe0f426bb2a8e7e,
	64'hbfe0f426bb2a8e7e, 64'h3feb23cd470013b4,
	64'h3fcccf8cb312b286, 64'h3fef2dc9c9089a9d,
	64'hbfef2dc9c9089a9d, 64'h3fcccf8cb312b286,
	64'h3feded05f7de47da, 64'h3fd6aa9d7dc77e17,
	64'hbfd6aa9d7dc77e17, 64'h3feded05f7de47da,
	64'h3fda4b4127dea1e5, 64'h3fed2cb220e0ef9f,
	64'hbfed2cb220e0ef9f, 64'h3fda4b4127dea1e5,
	64'h3fe74f948da8d28d, 64'h3fe5ec3495837074,
	64'hbfe5ec3495837074, 64'h3fe74f948da8d28d,
	64'h3f9f693731d1cf01, 64'h3feffc251df1d3f8,
	64'hbfeffc251df1d3f8, 64'h3f9f693731d1cf01,
	64'h3feff871dadb81df, 64'h3fa5fc00d290cd43,
	64'hbfa5fc00d290cd43, 64'h3feff871dadb81df,
	64'h3fe5a28d2a5d7250, 64'h3fe79400574f55e5,
	64'hbfe79400574f55e5, 64'h3fe5a28d2a5d7250,
	64'h3fed02d4feb2bd92, 64'h3fdb020d6c7f4009,
	64'hbfdb020d6c7f4009, 64'h3fed02d4feb2bd92,
	64'h3fd5ee27379ea693, 64'h3fee100cca2980ac,
	64'hbfee100cca2980ac, 64'h3fd5ee27379ea693,
	64'h3fef168f53f7205d, 64'h3fce56ca1e101a1b,
	64'hbfce56ca1e101a1b, 64'h3fef168f53f7205d,
	64'h3fe09e907417c5e1, 64'h3feb5889fe921405,
	64'hbfeb5889fe921405, 64'h3fe09e907417c5e1,
	64'h3fe9d1b1f5ea80d5, 64'h3fe2e780e3e8ea17,
	64'hbfe2e780e3e8ea17, 64'h3fe9d1b1f5ea80d5,
	64'h3fc38edbb0cd8d14, 64'h3fef9fce55adb2c8,
	64'hbfef9fce55adb2c8, 64'h3fc38edbb0cd8d14,
	64'h3fefae8e8e46cfbb, 64'h3fc20116d4ec7bcf,
	64'hbfc20116d4ec7bcf, 64'h3fefae8e8e46cfbb,
	64'h3fe338400d0c8e57, 64'h3fe995cf2ed80d22,
	64'hbfe995cf2ed80d22, 64'h3fe338400d0c8e57,
	64'h3feb8c38d27504e9, 64'h3fe0485626ae221a,
	64'hbfe0485626ae221a, 64'h3feb8c38d27504e9,
	64'h3fcfdcdc1adfedf9, 64'h3feefe220c0b95ec,
	64'hbfeefe220c0b95ec, 64'h3fcfdcdc1adfedf9,
	64'h3fee31eae870ce25, 64'h3fd530d880af3c24,
	64'hbfd530d880af3c24, 64'h3fee31eae870ce25,
	64'h3fdbb7cf2304bd01, 64'h3fecd7d9898b32f6,
	64'hbfecd7d9898b32f6, 64'h3fdbb7cf2304bd01,
	64'h3fe7d7836cc33db2, 64'h3fe5581038975137,
	64'hbfe5581038975137, 64'h3fe7d7836cc33db2,
	64'h3fac428d12c0d7e3, 64'h3feff3830f8d575c,
	64'hbfeff3830f8d575c, 64'h3fac428d12c0d7e3,
	64'h3fefdd539ff1f456, 64'h3fb787586a5d5b21,
	64'hbfb787586a5d5b21, 64'h3fefdd539ff1f456,
	64'h3fe473b51b987347, 64'h3fe89c7e9a4dd4aa,
	64'hbfe89c7e9a4dd4aa, 64'h3fe473b51b987347,
	64'h3fec5042012b6907, 64'h3fddd28f1481cc58,
	64'hbfddd28f1481cc58, 64'h3fec5042012b6907,
	64'h3fd2f422daec0387, 64'h3fee9084361df7f2,
	64'hbfee9084361df7f2, 64'h3fd2f422daec0387,
	64'h3feeadb2e8e7a88e, 64'h3fd233bbabc3bb71,
	64'hbfd233bbabc3bb71, 64'h3feeadb2e8e7a88e,
	64'h3fde83e0eaf85114, 64'h3fec20de3fa971b0,
	64'hbfec20de3fa971b0, 64'h3fde83e0eaf85114,
	64'h3fe8dc45331698cc, 64'h3fe425ff178e6bb1,
	64'hbfe425ff178e6bb1, 64'h3fe8dc45331698cc,
	64'h3fbaa7b724495c03, 64'h3fefd37914220b84,
	64'hbfefd37914220b84, 64'h3fbaa7b724495c03,
	64'h3fef6c3f7df5bbb7, 64'h3fc83366e89c64c6,
	64'hbfc83366e89c64c6, 64'h3fef6c3f7df5bbb7,
	64'h3fe1f0f08bbc861b, 64'h3fea7f58529fe69d,
	64'hbfea7f58529fe69d, 64'h3fe1f0f08bbc861b,
	64'h3feab7325916c0d4, 64'h3fe19d5a09f2b9b8,
	64'hbfe19d5a09f2b9b8, 64'h3feab7325916c0d4,
	64'h3fc9bdcbf2dc4366, 64'h3fef58a2b1789e84,
	64'hbfef58a2b1789e84, 64'h3fc9bdcbf2dc4366,
	64'h3feda383a9668988, 64'h3fd820e3b04eaac4,
	64'hbfd820e3b04eaac4, 64'h3feda383a9668988,
	64'h3fd8daa52ec8a4b0, 64'h3fed7d0b02b8ecf9,
	64'hbfed7d0b02b8ecf9, 64'h3fd8daa52ec8a4b0,
	64'h3fe6c40d73c18275, 64'h3fe67cf78491af10,
	64'hbfe67cf78491af10, 64'h3fe6c40d73c18275,
	64'h3f7921f0fe670071, 64'h3fefffd8858e8a92,
	64'hbfefffd8858e8a92, 64'h3f7921f0fe670071,
	64'h3feffff621621d02, 64'h3f6921f8becca4ba,
	64'hbf6921f8becca4ba, 64'h3feffff621621d02,
	64'h3fe68ed1eaa19c71, 64'h3fe6b25ced2fe29c,
	64'hbfe6b25ced2fe29c, 64'h3fe68ed1eaa19c71,
	64'h3fed86c48445a44f, 64'h3fd8ac4b86d5ed44,
	64'hbfd8ac4b86d5ed44, 64'h3fed86c48445a44f,
	64'h3fd84f6aaaf3903f, 64'h3fed9a00dd8b3d46,
	64'hbfed9a00dd8b3d46, 64'h3fd84f6aaaf3903f,
	64'h3fef5da6ed43685d, 64'h3fc95b49e9b62afa,
	64'hbfc95b49e9b62afa, 64'h3fef5da6ed43685d,
	64'h3fe1b250171373bf, 64'h3feaa9547a2cb98e,
	64'hbfeaa9547a2cb98e, 64'h3fe1b250171373bf,
	64'h3fea8d676e545ad2, 64'h3fe1dc1b64dc4872,
	64'hbfe1dc1b64dc4872, 64'h3fea8d676e545ad2,
	64'h3fc8961727c41804, 64'h3fef677556883cee,
	64'hbfef677556883cee, 64'h3fc8961727c41804,
	64'h3fefd60d2da75c9e, 64'h3fb9dfb6eb24a85c,
	64'hbfb9dfb6eb24a85c, 64'h3fefd60d2da75c9e,
	64'h3fe4397f5b2a4380, 64'h3fe8cc6a75184655,
	64'hbfe8cc6a75184655, 64'h3fe4397f5b2a4380,
	64'h3fec2cd14931e3f1, 64'h3fde57a86d3cd825,
	64'hbfde57a86d3cd825, 64'h3fec2cd14931e3f1,
	64'h3fd263e6995554ba, 64'h3feea68393e65800,
	64'hbfeea68393e65800, 64'h3fd263e6995554ba,
	64'h3fee97ec36016b30, 64'h3fd2c41a4e954520,
	64'hbfd2c41a4e954520, 64'h3fee97ec36016b30,
	64'h3fddfeff66a941de, 64'h3fec44833141c004,
	64'hbfec44833141c004, 64'h3fddfeff66a941de,
	64'h3fe8ac871ede1d88, 64'h3fe4605a692b32a2,
	64'hbfe4605a692b32a2, 64'h3fe8ac871ede1d88,
	64'h3fb84f8712c130a1, 64'h3fefdafa7514538c,
	64'hbfefdafa7514538c, 64'h3fb84f8712c130a1,
	64'h3feff4dc54b1bed3, 64'h3faab101bd5f8317,
	64'hbfaab101bd5f8317, 64'h3feff4dc54b1bed3,
	64'h3fe56ac35197649f, 64'h3fe7c6b89ce2d333,
	64'hbfe7c6b89ce2d333, 64'h3fe56ac35197649f,
	64'h3fece2b32799a060, 64'h3fdb8a7814fd5693,
	64'hbfdb8a7814fd5693, 64'h3fece2b32799a060,
	64'h3fd5604012f467b4, 64'h3fee298f4439197a,
	64'hbfee298f4439197a, 64'h3fd5604012f467b4,
	64'h3fef045a14cf738c, 64'h3fcf7b7480bd3802,
	64'hbfcf7b7480bd3802, 64'h3fef045a14cf738c,
	64'h3fe05df3ec31b8b7, 64'h3feb7f6686e792e9,
	64'hbfeb7f6686e792e9, 64'h3fe05df3ec31b8b7,
	64'h3fe9a4dfa42b06b2, 64'h3fe32421ec49a61f,
	64'hbfe32421ec49a61f, 64'h3fe9a4dfa42b06b2,
	64'h3fc264994dfd3409, 64'h3fefaafbcb0cfddc,
	64'hbfefaafbcb0cfddc, 64'h3fc264994dfd3409,
	64'h3fefa39bac7a1791, 64'h3fc32b7bf94516a7,
	64'hbfc32b7bf94516a7, 64'h3fefa39bac7a1791,
	64'h3fe2fbc24b441015, 64'h3fe9c2d110f075c2,
	64'hbfe9c2d110f075c2, 64'h3fe2fbc24b441015,
	64'h3feb658f14fdbc47, 64'h3fe089112032b08c,
	64'hbfe089112032b08c, 64'h3feb658f14fdbc47,
	64'h3fceb86b462de348, 64'h3fef1090bc898f5f,
	64'hbfef1090bc898f5f, 64'h3fceb86b462de348,
	64'h3fee18a02fdc66d9, 64'h3fd5bee78b9db3b6,
	64'hbfd5bee78b9db3b6, 64'h3fee18a02fdc66d9,
	64'h3fdb2f971db31972, 64'h3fecf830e8ce467b,
	64'hbfecf830e8ce467b, 64'h3fdb2f971db31972,
	64'h3fe7a4f707bf97d2, 64'h3fe59001d5f723df,
	64'hbfe59001d5f723df, 64'h3fe7a4f707bf97d2,
	64'h3fa78dbaa5874686, 64'h3feff753bb1b9164,
	64'hbfeff753bb1b9164, 64'h3fa78dbaa5874686,
	64'h3feffce09ce2a679, 64'h3f9c454f4ce53b1d,
	64'hbf9c454f4ce53b1d, 64'h3feffce09ce2a679,
	64'h3fe5fe7cbde56a10, 64'h3fe73e558e079942,
	64'hbfe73e558e079942, 64'h3fe5fe7cbde56a10,
	64'h3fed36fc7bcbfbdc, 64'h3fda1d6543b50ac0,
	64'hbfda1d6543b50ac0, 64'h3fed36fc7bcbfbdc,
	64'h3fd6d998638a0cb6, 64'h3fede4160f6d8d81,
	64'hbfede4160f6d8d81, 64'h3fd6d998638a0cb6,
	64'h3fef33685a3aaef0, 64'h3fcc6d90535d74dd,
	64'hbfcc6d90535d74dd, 64'h3fef33685a3aaef0,
	64'h3fe1097248d0a957, 64'h3feb16742a4ca2f5,
	64'hbfeb16742a4ca2f5, 64'h3fe1097248d0a957,
	64'h3fea1b26d2c0a75e, 64'h3fe2818bef4d3cba,
	64'hbfe2818bef4d3cba, 64'h3fea1b26d2c0a75e,
	64'h3fc57f008654cbde, 64'h3fef8ba737cb4b78,
	64'hbfef8ba737cb4b78, 64'h3fc57f008654cbde,
	64'h3fefbf470f0a8d88, 64'h3fc00ee8ad6fb85b,
	64'hbfc00ee8ad6fb85b, 64'h3fefbf470f0a8d88,
	64'h3fe39c23e3d63029, 64'h3fe94990e3ac4a6c,
	64'hbfe94990e3ac4a6c, 64'h3fe39c23e3d63029,
	64'h3febcb54cb0d2327, 64'h3fdfb7575c24d2de,
	64'hbfdfb7575c24d2de, 64'h3febcb54cb0d2327,
	64'h3fd0e15b4e1749ce, 64'h3feeddeb6a078651,
	64'hbfeeddeb6a078651, 64'h3fd0e15b4e1749ce,
	64'h3fee5a9d550467d3, 64'h3fd44310dc8936f0,
	64'hbfd44310dc8936f0, 64'h3fee5a9d550467d3,
	64'h3fdc997fc3865389, 64'h3feca08f19b9c449,
	64'hbfeca08f19b9c449, 64'h3fdc997fc3865389,
	64'h3fe82a9c13f545ff, 64'h3fe4f9cc25cca486,
	64'hbfe4f9cc25cca486, 64'h3fe82a9c13f545ff,
	64'h3fb20c9674ed444d, 64'h3fefeb9d2530410f,
	64'hbfefeb9d2530410f, 64'h3fb20c9674ed444d,
	64'h3fefe7ea85482d60, 64'h3fb39d9f12c5a299,
	64'hbfb39d9f12c5a299, 64'h3fefe7ea85482d60,
	64'h3fe4d3bc6d589f7f, 64'h3fe84b7111af83fa,
	64'hbfe84b7111af83fa, 64'h3fe4d3bc6d589f7f,
	64'h3fec89f587029c13, 64'h3fdcf34baee1cd21,
	64'hbfdcf34baee1cd21, 64'h3fec89f587029c13,
	64'h3fd3e39be96ec271, 64'h3fee6a61c55d53a7,
	64'hbfee6a61c55d53a7, 64'h3fd3e39be96ec271,
	64'h3feed0835e999009, 64'h3fd1423eefc69378,
	64'hbfd1423eefc69378, 64'h3feed0835e999009,
	64'h3fdf5fdee656cda3, 64'h3febe41b611154c1,
	64'hbfebe41b611154c1, 64'h3fdf5fdee656cda3,
	64'h3fe92aa41fc5a815, 64'h3fe3c3c44981c518,
	64'hbfe3c3c44981c518, 64'h3fe92aa41fc5a815,
	64'h3fbe8eb7fde4aa3f, 64'h3fefc56e3b7d9af6,
	64'hbfefc56e3b7d9af6, 64'h3fbe8eb7fde4aa3f,
	64'h3fef830f4a40c60c, 64'h3fc6451a831d830d,
	64'hbfc6451a831d830d, 64'h3fef830f4a40c60c,
	64'h3fe258734cbb7110, 64'h3fea38184a593bc6,
	64'hbfea38184a593bc6, 64'h3fe258734cbb7110,
	64'h3feafb8fd89f57b6, 64'h3fe133e9cfee254f,
	64'hbfe133e9cfee254f, 64'h3feafb8fd89f57b6,
	64'h3fcba96334f15dad, 64'h3fef3e6bbc1bbc65,
	64'hbfef3e6bbc1bbc65, 64'h3fcba96334f15dad,
	64'h3fedd1fef38a915a, 64'h3fd73763c9261092,
	64'hbfd73763c9261092, 64'h3fedd1fef38a915a,
	64'h3fd9c17d440df9f2, 64'h3fed4b5b1b187524,
	64'hbfed4b5b1b187524, 64'h3fd9c17d440df9f2,
	64'h3fe71bac960e41bf, 64'h3fe622e44fec22ff,
	64'hbfe622e44fec22ff, 64'h3fe71bac960e41bf,
	64'h3f95fd4d21fab226, 64'h3feffe1c6870cb77,
	64'hbfeffe1c6870cb77, 64'h3f95fd4d21fab226,
	64'h3fefff0943c53bd1, 64'h3f8f6a296ab997cb,
	64'hbf8f6a296ab997cb, 64'h3fefff0943c53bd1,
	64'h3fe64715437f535b, 64'h3fe6f8ca99c95b75,
	64'hbfe6f8ca99c95b75, 64'h3fe64715437f535b,
	64'h3fed5f7172888a7f, 64'h3fd96555b7ab948f,
	64'hbfd96555b7ab948f, 64'h3fed5f7172888a7f,
	64'h3fd794f5e613dfae, 64'h3fedbf9e4395759a,
	64'hbfedbf9e4395759a, 64'h3fd794f5e613dfae,
	64'h3fef492206bcabb4, 64'h3fcae4f1d5f3b9ab,
	64'hbfcae4f1d5f3b9ab, 64'h3fef492206bcabb4,
	64'h3fe15e36e4dbe2bc, 64'h3feae068f345ecef,
	64'hbfeae068f345ecef, 64'h3fe15e36e4dbe2bc,
	64'h3fea54c91090f523, 64'h3fe22f2d662c13e2,
	64'hbfe22f2d662c13e2, 64'h3fea54c91090f523,
	64'h3fc70afd8d08c4ff, 64'h3fef7a299c1a322a,
	64'hbfef7a299c1a322a, 64'h3fc70afd8d08c4ff,
	64'h3fefcb4703914354, 64'h3fbcff533b307dc1,
	64'hbfbcff533b307dc1, 64'h3fefcb4703914354,
	64'h3fe3eb33eabe0680, 64'h3fe90b7943575efe,
	64'hbfe90b7943575efe, 64'h3fe3eb33eabe0680,
	64'h3febfc9d25a1b147, 64'h3fdf081906bff7fe,
	64'hbfdf081906bff7fe, 64'h3febfc9d25a1b147,
	64'h3fd1a2f7fbe8f243, 64'h3feec2cf4b1af6b2,
	64'hbfeec2cf4b1af6b2, 64'h3fd1a2f7fbe8f243,
	64'h3fee79db29a5165a, 64'h3fd383f5e353b6ab,
	64'hbfd383f5e353b6ab, 64'h3fee79db29a5165a,
	64'h3fdd4cd02ba8609d, 64'h3fec7315899eaad7,
	64'hbfec7315899eaad7, 64'h3fdd4cd02ba8609d,
	64'h3fe86c0a1d9aa195, 64'h3fe4ad79516722f1,
	64'hbfe4ad79516722f1, 64'h3fe86c0a1d9aa195,
	64'h3fb52e774a4d4d0a, 64'h3fefe3e92be9d886,
	64'hbfefe3e92be9d886, 64'h3fb52e774a4d4d0a,
	64'h3fefef0102826191, 64'h3fb07b614e463064,
	64'hbfb07b614e463064, 64'h3fefef0102826191,
	64'h3fe51fa81cd99aa6, 64'h3fe8098b756e52fa,
	64'hbfe8098b756e52fa, 64'h3fe51fa81cd99aa6,
	64'h3fecb6e20a00da99, 64'h3fdc3f6d47263129,
	64'hbfdc3f6d47263129, 64'h3fecb6e20a00da99,
	64'h3fd4a253d11b82f3, 64'h3fee4a8dff81ce5e,
	64'hbfee4a8dff81ce5e, 64'h3fd4a253d11b82f3,
	64'h3feeeb074c50a544, 64'h3fd0804e05eb661e,
	64'hbfd0804e05eb661e, 64'h3feeeb074c50a544,
	64'h3fe00740c82b82e1, 64'h3febb249a0b6c40d,
	64'hbfebb249a0b6c40d, 64'h3fe00740c82b82e1,
	64'h3fe9683f42bd7fe1, 64'h3fe374531b817f8d,
	64'hbfe374531b817f8d, 64'h3fe9683f42bd7fe1,
	64'h3fc0d64dbcb26786, 64'h3fefb8d18d66adb7,
	64'hbfefb8d18d66adb7, 64'h3fc0d64dbcb26786,
	64'h3fef93f14f85ac08, 64'h3fc4b8b17f79fa88,
	64'hbfc4b8b17f79fa88, 64'h3fef93f14f85ac08,
	64'h3fe2aa76e87aeb58, 64'h3fe9fdf4f13149de,
	64'hbfe9fdf4f13149de, 64'h3fe2aa76e87aeb58,
	64'h3feb3115a5f37bf3, 64'h3fe0ded0b84bc4b6,
	64'hbfe0ded0b84bc4b6, 64'h3feb3115a5f37bf3,
	64'h3fcd31774d2cbdee, 64'h3fef2817fc4609ce,
	64'hbfef2817fc4609ce, 64'h3fcd31774d2cbdee,
	64'h3fedf5e36a9ba59c, 64'h3fd67b949cad63cb,
	64'hbfd67b949cad63cb, 64'h3fedf5e36a9ba59c,
	64'h3fda790cd3dbf31b, 64'h3fed2255c6e5a4e1,
	64'hbfed2255c6e5a4e1, 64'h3fda790cd3dbf31b,
	64'h3fe760c52c304764, 64'h3fe5d9dee73e345c,
	64'hbfe5d9dee73e345c, 64'h3fe760c52c304764,
	64'h3fa14685db42c17f, 64'h3feffb55e425fdae,
	64'hbfeffb55e425fdae, 64'h3fa14685db42c17f,
	64'h3feff97c4208c014, 64'h3fa46a396ff86179,
	64'hbfa46a396ff86179, 64'h3feff97c4208c014,
	64'h3fe5b50b264f7448, 64'h3fe782fb1b90b35b,
	64'hbfe782fb1b90b35b, 64'h3fe5b50b264f7448,
	64'h3fed0d672f59d2b9, 64'h3fdad473125cdc09,
	64'hbfdad473125cdc09, 64'h3fed0d672f59d2b9,
	64'h3fd61d595c88c202, 64'h3fee0766d9280f54,
	64'hbfee0766d9280f54, 64'h3fd61d595c88c202,
	64'h3fef1c7abe284708, 64'h3fcdf5163f01099a,
	64'hbfcdf5163f01099a, 64'h3fef1c7abe284708,
	64'h3fe0b405878f85ec, 64'h3feb4b7409de7925,
	64'hbfeb4b7409de7925, 64'h3fe0b405878f85ec,
	64'h3fe9e082edb42472, 64'h3fe2d333d34e9bb8,
	64'hbfe2d333d34e9bb8, 64'h3fe9e082edb42472,
	64'h3fc3f22f57db4893, 64'h3fef9bed7cfbde29,
	64'hbfef9bed7cfbde29, 64'h3fc3f22f57db4893,
	64'h3fefb20dc681d54d, 64'h3fc19d8940be24e7,
	64'hbfc19d8940be24e7, 64'h3fefb20dc681d54d,
	64'h3fe34c5252c14de1, 64'h3fe986aef1457594,
	64'hbfe986aef1457594, 64'h3fe34c5252c14de1,
	64'h3feb98fa1fd9155e, 64'h3fe032ae55edbd96,
	64'hbfe032ae55edbd96, 64'h3feb98fa1fd9155e,
	64'h3fd01f1806b9fdd2, 64'h3feef7d6e51ca3c0,
	64'hbfeef7d6e51ca3c0, 64'h3fd01f1806b9fdd2,
	64'h3fee3a33ec75ce85, 64'h3fd50163dc197048,
	64'hbfd50163dc197048, 64'h3fee3a33ec75ce85,
	64'h3fdbe51517ffc0d9, 64'h3fecccee20c2dea0,
	64'hbfecccee20c2dea0, 64'h3fdbe51517ffc0d9,
	64'h3fe7e83f87b03686, 64'h3fe5454ff5159dfc,
	64'hbfe5454ff5159dfc, 64'h3fe7e83f87b03686,
	64'h3fadd406f9808ec9, 64'h3feff21614e131ed,
	64'hbfeff21614e131ed, 64'h3fadd406f9808ec9,
	64'h3fefdf9922f73307, 64'h3fb6bf1b3e79b129,
	64'hbfb6bf1b3e79b129, 64'h3fefdf9922f73307,
	64'h3fe48703306091ff, 64'h3fe88c66e7481ba1,
	64'hbfe88c66e7481ba1, 64'h3fe48703306091ff,
	64'h3fec5bef59fef85a, 64'h3fdda60c5cfa10d9,
	64'hbfdda60c5cfa10d9, 64'h3fec5bef59fef85a,
	64'h3fd3241fb638baaf, 64'h3fee89095bad6025,
	64'hbfee89095bad6025, 64'h3fd3241fb638baaf,
	64'h3feeb4cf515b8811, 64'h3fd2038583d727be,
	64'hbfd2038583d727be, 64'h3feeb4cf515b8811,
	64'h3fdeb00695f25620, 64'h3fec14d9dc465e57,
	64'hbfec14d9dc465e57, 64'h3fdeb00695f25620,
	64'h3fe8ec109b486c49, 64'h3fe41272663d108c,
	64'hbfe41272663d108c, 64'h3fe8ec109b486c49,
	64'h3fbb6fa6ec38f64c, 64'h3fefd0d158d86087,
	64'hbfefd0d158d86087, 64'h3fbb6fa6ec38f64c,
	64'h3fef70f6434b7eb7, 64'h3fc7d0a7bbd2cb1c,
	64'hbfc7d0a7bbd2cb1c, 64'h3fef70f6434b7eb7,
	64'h3fe205baa17560d6, 64'h3fea7138de9d60f5,
	64'hbfea7138de9d60f5, 64'h3fe205baa17560d6,
	64'h3feac4ffbd3efac8, 64'h3fe188591f3a46e5,
	64'hbfe188591f3a46e5, 64'h3feac4ffbd3efac8,
	64'h3fca203e1b1831da, 64'h3fef538b1faf2d07,
	64'hbfef538b1faf2d07, 64'h3fca203e1b1831da,
	64'h3fedacf42ce68ab9, 64'h3fd7f24dd37341e4,
	64'hbfd7f24dd37341e4, 64'h3fedacf42ce68ab9,
	64'h3fd908ef81ef7bd1, 64'h3fed733f508c0dff,
	64'hbfed733f508c0dff, 64'h3fd908ef81ef7bd1,
	64'h3fe6d5afef4aafcd, 64'h3fe66b0f3f52b386,
	64'hbfe66b0f3f52b386, 64'h3fe6d5afef4aafcd,
	64'h3f82d96b0e509703, 64'h3fefffa72c978c4f,
	64'hbfefffa72c978c4f, 64'h3f82d96b0e509703,
	64'h3fefffa72c978c4f, 64'h3f82d96b0e509703,
	64'hbf82d96b0e509703, 64'h3fefffa72c978c4f,
	64'h3fe66b0f3f52b386, 64'h3fe6d5afef4aafcd,
	64'hbfe6d5afef4aafcd, 64'h3fe66b0f3f52b386,
	64'h3fed733f508c0dff, 64'h3fd908ef81ef7bd1,
	64'hbfd908ef81ef7bd1, 64'h3fed733f508c0dff,
	64'h3fd7f24dd37341e4, 64'h3fedacf42ce68ab9,
	64'hbfedacf42ce68ab9, 64'h3fd7f24dd37341e4,
	64'h3fef538b1faf2d07, 64'h3fca203e1b1831da,
	64'hbfca203e1b1831da, 64'h3fef538b1faf2d07,
	64'h3fe188591f3a46e5, 64'h3feac4ffbd3efac8,
	64'hbfeac4ffbd3efac8, 64'h3fe188591f3a46e5,
	64'h3fea7138de9d60f5, 64'h3fe205baa17560d6,
	64'hbfe205baa17560d6, 64'h3fea7138de9d60f5,
	64'h3fc7d0a7bbd2cb1c, 64'h3fef70f6434b7eb7,
	64'hbfef70f6434b7eb7, 64'h3fc7d0a7bbd2cb1c,
	64'h3fefd0d158d86087, 64'h3fbb6fa6ec38f64c,
	64'hbfbb6fa6ec38f64c, 64'h3fefd0d158d86087,
	64'h3fe41272663d108c, 64'h3fe8ec109b486c49,
	64'hbfe8ec109b486c49, 64'h3fe41272663d108c,
	64'h3fec14d9dc465e57, 64'h3fdeb00695f25620,
	64'hbfdeb00695f25620, 64'h3fec14d9dc465e57,
	64'h3fd2038583d727be, 64'h3feeb4cf515b8811,
	64'hbfeeb4cf515b8811, 64'h3fd2038583d727be,
	64'h3fee89095bad6025, 64'h3fd3241fb638baaf,
	64'hbfd3241fb638baaf, 64'h3fee89095bad6025,
	64'h3fdda60c5cfa10d9, 64'h3fec5bef59fef85a,
	64'hbfec5bef59fef85a, 64'h3fdda60c5cfa10d9,
	64'h3fe88c66e7481ba1, 64'h3fe48703306091ff,
	64'hbfe48703306091ff, 64'h3fe88c66e7481ba1,
	64'h3fb6bf1b3e79b129, 64'h3fefdf9922f73307,
	64'hbfefdf9922f73307, 64'h3fb6bf1b3e79b129,
	64'h3feff21614e131ed, 64'h3fadd406f9808ec9,
	64'hbfadd406f9808ec9, 64'h3feff21614e131ed,
	64'h3fe5454ff5159dfc, 64'h3fe7e83f87b03686,
	64'hbfe7e83f87b03686, 64'h3fe5454ff5159dfc,
	64'h3fecccee20c2dea0, 64'h3fdbe51517ffc0d9,
	64'hbfdbe51517ffc0d9, 64'h3fecccee20c2dea0,
	64'h3fd50163dc197048, 64'h3fee3a33ec75ce85,
	64'hbfee3a33ec75ce85, 64'h3fd50163dc197048,
	64'h3feef7d6e51ca3c0, 64'h3fd01f1806b9fdd2,
	64'hbfd01f1806b9fdd2, 64'h3feef7d6e51ca3c0,
	64'h3fe032ae55edbd96, 64'h3feb98fa1fd9155e,
	64'hbfeb98fa1fd9155e, 64'h3fe032ae55edbd96,
	64'h3fe986aef1457594, 64'h3fe34c5252c14de1,
	64'hbfe34c5252c14de1, 64'h3fe986aef1457594,
	64'h3fc19d8940be24e7, 64'h3fefb20dc681d54d,
	64'hbfefb20dc681d54d, 64'h3fc19d8940be24e7,
	64'h3fef9bed7cfbde29, 64'h3fc3f22f57db4893,
	64'hbfc3f22f57db4893, 64'h3fef9bed7cfbde29,
	64'h3fe2d333d34e9bb8, 64'h3fe9e082edb42472,
	64'hbfe9e082edb42472, 64'h3fe2d333d34e9bb8,
	64'h3feb4b7409de7925, 64'h3fe0b405878f85ec,
	64'hbfe0b405878f85ec, 64'h3feb4b7409de7925,
	64'h3fcdf5163f01099a, 64'h3fef1c7abe284708,
	64'hbfef1c7abe284708, 64'h3fcdf5163f01099a,
	64'h3fee0766d9280f54, 64'h3fd61d595c88c202,
	64'hbfd61d595c88c202, 64'h3fee0766d9280f54,
	64'h3fdad473125cdc09, 64'h3fed0d672f59d2b9,
	64'hbfed0d672f59d2b9, 64'h3fdad473125cdc09,
	64'h3fe782fb1b90b35b, 64'h3fe5b50b264f7448,
	64'hbfe5b50b264f7448, 64'h3fe782fb1b90b35b,
	64'h3fa46a396ff86179, 64'h3feff97c4208c014,
	64'hbfeff97c4208c014, 64'h3fa46a396ff86179,
	64'h3feffb55e425fdae, 64'h3fa14685db42c17f,
	64'hbfa14685db42c17f, 64'h3feffb55e425fdae,
	64'h3fe5d9dee73e345c, 64'h3fe760c52c304764,
	64'hbfe760c52c304764, 64'h3fe5d9dee73e345c,
	64'h3fed2255c6e5a4e1, 64'h3fda790cd3dbf31b,
	64'hbfda790cd3dbf31b, 64'h3fed2255c6e5a4e1,
	64'h3fd67b949cad63cb, 64'h3fedf5e36a9ba59c,
	64'hbfedf5e36a9ba59c, 64'h3fd67b949cad63cb,
	64'h3fef2817fc4609ce, 64'h3fcd31774d2cbdee,
	64'hbfcd31774d2cbdee, 64'h3fef2817fc4609ce,
	64'h3fe0ded0b84bc4b6, 64'h3feb3115a5f37bf3,
	64'hbfeb3115a5f37bf3, 64'h3fe0ded0b84bc4b6,
	64'h3fe9fdf4f13149de, 64'h3fe2aa76e87aeb58,
	64'hbfe2aa76e87aeb58, 64'h3fe9fdf4f13149de,
	64'h3fc4b8b17f79fa88, 64'h3fef93f14f85ac08,
	64'hbfef93f14f85ac08, 64'h3fc4b8b17f79fa88,
	64'h3fefb8d18d66adb7, 64'h3fc0d64dbcb26786,
	64'hbfc0d64dbcb26786, 64'h3fefb8d18d66adb7,
	64'h3fe374531b817f8d, 64'h3fe9683f42bd7fe1,
	64'hbfe9683f42bd7fe1, 64'h3fe374531b817f8d,
	64'h3febb249a0b6c40d, 64'h3fe00740c82b82e1,
	64'hbfe00740c82b82e1, 64'h3febb249a0b6c40d,
	64'h3fd0804e05eb661e, 64'h3feeeb074c50a544,
	64'hbfeeeb074c50a544, 64'h3fd0804e05eb661e,
	64'h3fee4a8dff81ce5e, 64'h3fd4a253d11b82f3,
	64'hbfd4a253d11b82f3, 64'h3fee4a8dff81ce5e,
	64'h3fdc3f6d47263129, 64'h3fecb6e20a00da99,
	64'hbfecb6e20a00da99, 64'h3fdc3f6d47263129,
	64'h3fe8098b756e52fa, 64'h3fe51fa81cd99aa6,
	64'hbfe51fa81cd99aa6, 64'h3fe8098b756e52fa,
	64'h3fb07b614e463064, 64'h3fefef0102826191,
	64'hbfefef0102826191, 64'h3fb07b614e463064,
	64'h3fefe3e92be9d886, 64'h3fb52e774a4d4d0a,
	64'hbfb52e774a4d4d0a, 64'h3fefe3e92be9d886,
	64'h3fe4ad79516722f1, 64'h3fe86c0a1d9aa195,
	64'hbfe86c0a1d9aa195, 64'h3fe4ad79516722f1,
	64'h3fec7315899eaad7, 64'h3fdd4cd02ba8609d,
	64'hbfdd4cd02ba8609d, 64'h3fec7315899eaad7,
	64'h3fd383f5e353b6ab, 64'h3fee79db29a5165a,
	64'hbfee79db29a5165a, 64'h3fd383f5e353b6ab,
	64'h3feec2cf4b1af6b2, 64'h3fd1a2f7fbe8f243,
	64'hbfd1a2f7fbe8f243, 64'h3feec2cf4b1af6b2,
	64'h3fdf081906bff7fe, 64'h3febfc9d25a1b147,
	64'hbfebfc9d25a1b147, 64'h3fdf081906bff7fe,
	64'h3fe90b7943575efe, 64'h3fe3eb33eabe0680,
	64'hbfe3eb33eabe0680, 64'h3fe90b7943575efe,
	64'h3fbcff533b307dc1, 64'h3fefcb4703914354,
	64'hbfefcb4703914354, 64'h3fbcff533b307dc1,
	64'h3fef7a299c1a322a, 64'h3fc70afd8d08c4ff,
	64'hbfc70afd8d08c4ff, 64'h3fef7a299c1a322a,
	64'h3fe22f2d662c13e2, 64'h3fea54c91090f523,
	64'hbfea54c91090f523, 64'h3fe22f2d662c13e2,
	64'h3feae068f345ecef, 64'h3fe15e36e4dbe2bc,
	64'hbfe15e36e4dbe2bc, 64'h3feae068f345ecef,
	64'h3fcae4f1d5f3b9ab, 64'h3fef492206bcabb4,
	64'hbfef492206bcabb4, 64'h3fcae4f1d5f3b9ab,
	64'h3fedbf9e4395759a, 64'h3fd794f5e613dfae,
	64'hbfd794f5e613dfae, 64'h3fedbf9e4395759a,
	64'h3fd96555b7ab948f, 64'h3fed5f7172888a7f,
	64'hbfed5f7172888a7f, 64'h3fd96555b7ab948f,
	64'h3fe6f8ca99c95b75, 64'h3fe64715437f535b,
	64'hbfe64715437f535b, 64'h3fe6f8ca99c95b75,
	64'h3f8f6a296ab997cb, 64'h3fefff0943c53bd1,
	64'hbfefff0943c53bd1, 64'h3f8f6a296ab997cb,
	64'h3feffe1c6870cb77, 64'h3f95fd4d21fab226,
	64'hbf95fd4d21fab226, 64'h3feffe1c6870cb77,
	64'h3fe622e44fec22ff, 64'h3fe71bac960e41bf,
	64'hbfe71bac960e41bf, 64'h3fe622e44fec22ff,
	64'h3fed4b5b1b187524, 64'h3fd9c17d440df9f2,
	64'hbfd9c17d440df9f2, 64'h3fed4b5b1b187524,
	64'h3fd73763c9261092, 64'h3fedd1fef38a915a,
	64'hbfedd1fef38a915a, 64'h3fd73763c9261092,
	64'h3fef3e6bbc1bbc65, 64'h3fcba96334f15dad,
	64'hbfcba96334f15dad, 64'h3fef3e6bbc1bbc65,
	64'h3fe133e9cfee254f, 64'h3feafb8fd89f57b6,
	64'hbfeafb8fd89f57b6, 64'h3fe133e9cfee254f,
	64'h3fea38184a593bc6, 64'h3fe258734cbb7110,
	64'hbfe258734cbb7110, 64'h3fea38184a593bc6,
	64'h3fc6451a831d830d, 64'h3fef830f4a40c60c,
	64'hbfef830f4a40c60c, 64'h3fc6451a831d830d,
	64'h3fefc56e3b7d9af6, 64'h3fbe8eb7fde4aa3f,
	64'hbfbe8eb7fde4aa3f, 64'h3fefc56e3b7d9af6,
	64'h3fe3c3c44981c518, 64'h3fe92aa41fc5a815,
	64'hbfe92aa41fc5a815, 64'h3fe3c3c44981c518,
	64'h3febe41b611154c1, 64'h3fdf5fdee656cda3,
	64'hbfdf5fdee656cda3, 64'h3febe41b611154c1,
	64'h3fd1423eefc69378, 64'h3feed0835e999009,
	64'hbfeed0835e999009, 64'h3fd1423eefc69378,
	64'h3fee6a61c55d53a7, 64'h3fd3e39be96ec271,
	64'hbfd3e39be96ec271, 64'h3fee6a61c55d53a7,
	64'h3fdcf34baee1cd21, 64'h3fec89f587029c13,
	64'hbfec89f587029c13, 64'h3fdcf34baee1cd21,
	64'h3fe84b7111af83fa, 64'h3fe4d3bc6d589f7f,
	64'hbfe4d3bc6d589f7f, 64'h3fe84b7111af83fa,
	64'h3fb39d9f12c5a299, 64'h3fefe7ea85482d60,
	64'hbfefe7ea85482d60, 64'h3fb39d9f12c5a299,
	64'h3fefeb9d2530410f, 64'h3fb20c9674ed444d,
	64'hbfb20c9674ed444d, 64'h3fefeb9d2530410f,
	64'h3fe4f9cc25cca486, 64'h3fe82a9c13f545ff,
	64'hbfe82a9c13f545ff, 64'h3fe4f9cc25cca486,
	64'h3feca08f19b9c449, 64'h3fdc997fc3865389,
	64'hbfdc997fc3865389, 64'h3feca08f19b9c449,
	64'h3fd44310dc8936f0, 64'h3fee5a9d550467d3,
	64'hbfee5a9d550467d3, 64'h3fd44310dc8936f0,
	64'h3feeddeb6a078651, 64'h3fd0e15b4e1749ce,
	64'hbfd0e15b4e1749ce, 64'h3feeddeb6a078651,
	64'h3fdfb7575c24d2de, 64'h3febcb54cb0d2327,
	64'hbfebcb54cb0d2327, 64'h3fdfb7575c24d2de,
	64'h3fe94990e3ac4a6c, 64'h3fe39c23e3d63029,
	64'hbfe39c23e3d63029, 64'h3fe94990e3ac4a6c,
	64'h3fc00ee8ad6fb85b, 64'h3fefbf470f0a8d88,
	64'hbfefbf470f0a8d88, 64'h3fc00ee8ad6fb85b,
	64'h3fef8ba737cb4b78, 64'h3fc57f008654cbde,
	64'hbfc57f008654cbde, 64'h3fef8ba737cb4b78,
	64'h3fe2818bef4d3cba, 64'h3fea1b26d2c0a75e,
	64'hbfea1b26d2c0a75e, 64'h3fe2818bef4d3cba,
	64'h3feb16742a4ca2f5, 64'h3fe1097248d0a957,
	64'hbfe1097248d0a957, 64'h3feb16742a4ca2f5,
	64'h3fcc6d90535d74dd, 64'h3fef33685a3aaef0,
	64'hbfef33685a3aaef0, 64'h3fcc6d90535d74dd,
	64'h3fede4160f6d8d81, 64'h3fd6d998638a0cb6,
	64'hbfd6d998638a0cb6, 64'h3fede4160f6d8d81,
	64'h3fda1d6543b50ac0, 64'h3fed36fc7bcbfbdc,
	64'hbfed36fc7bcbfbdc, 64'h3fda1d6543b50ac0,
	64'h3fe73e558e079942, 64'h3fe5fe7cbde56a10,
	64'hbfe5fe7cbde56a10, 64'h3fe73e558e079942,
	64'h3f9c454f4ce53b1d, 64'h3feffce09ce2a679,
	64'hbfeffce09ce2a679, 64'h3f9c454f4ce53b1d,
	64'h3feff753bb1b9164, 64'h3fa78dbaa5874686,
	64'hbfa78dbaa5874686, 64'h3feff753bb1b9164,
	64'h3fe59001d5f723df, 64'h3fe7a4f707bf97d2,
	64'hbfe7a4f707bf97d2, 64'h3fe59001d5f723df,
	64'h3fecf830e8ce467b, 64'h3fdb2f971db31972,
	64'hbfdb2f971db31972, 64'h3fecf830e8ce467b,
	64'h3fd5bee78b9db3b6, 64'h3fee18a02fdc66d9,
	64'hbfee18a02fdc66d9, 64'h3fd5bee78b9db3b6,
	64'h3fef1090bc898f5f, 64'h3fceb86b462de348,
	64'hbfceb86b462de348, 64'h3fef1090bc898f5f,
	64'h3fe089112032b08c, 64'h3feb658f14fdbc47,
	64'hbfeb658f14fdbc47, 64'h3fe089112032b08c,
	64'h3fe9c2d110f075c2, 64'h3fe2fbc24b441015,
	64'hbfe2fbc24b441015, 64'h3fe9c2d110f075c2,
	64'h3fc32b7bf94516a7, 64'h3fefa39bac7a1791,
	64'hbfefa39bac7a1791, 64'h3fc32b7bf94516a7,
	64'h3fefaafbcb0cfddc, 64'h3fc264994dfd3409,
	64'hbfc264994dfd3409, 64'h3fefaafbcb0cfddc,
	64'h3fe32421ec49a61f, 64'h3fe9a4dfa42b06b2,
	64'hbfe9a4dfa42b06b2, 64'h3fe32421ec49a61f,
	64'h3feb7f6686e792e9, 64'h3fe05df3ec31b8b7,
	64'hbfe05df3ec31b8b7, 64'h3feb7f6686e792e9,
	64'h3fcf7b7480bd3802, 64'h3fef045a14cf738c,
	64'hbfef045a14cf738c, 64'h3fcf7b7480bd3802,
	64'h3fee298f4439197a, 64'h3fd5604012f467b4,
	64'hbfd5604012f467b4, 64'h3fee298f4439197a,
	64'h3fdb8a7814fd5693, 64'h3fece2b32799a060,
	64'hbfece2b32799a060, 64'h3fdb8a7814fd5693,
	64'h3fe7c6b89ce2d333, 64'h3fe56ac35197649f,
	64'hbfe56ac35197649f, 64'h3fe7c6b89ce2d333,
	64'h3faab101bd5f8317, 64'h3feff4dc54b1bed3,
	64'hbfeff4dc54b1bed3, 64'h3faab101bd5f8317,
	64'h3fefdafa7514538c, 64'h3fb84f8712c130a1,
	64'hbfb84f8712c130a1, 64'h3fefdafa7514538c,
	64'h3fe4605a692b32a2, 64'h3fe8ac871ede1d88,
	64'hbfe8ac871ede1d88, 64'h3fe4605a692b32a2,
	64'h3fec44833141c004, 64'h3fddfeff66a941de,
	64'hbfddfeff66a941de, 64'h3fec44833141c004,
	64'h3fd2c41a4e954520, 64'h3fee97ec36016b30,
	64'hbfee97ec36016b30, 64'h3fd2c41a4e954520,
	64'h3feea68393e65800, 64'h3fd263e6995554ba,
	64'hbfd263e6995554ba, 64'h3feea68393e65800,
	64'h3fde57a86d3cd825, 64'h3fec2cd14931e3f1,
	64'hbfec2cd14931e3f1, 64'h3fde57a86d3cd825,
	64'h3fe8cc6a75184655, 64'h3fe4397f5b2a4380,
	64'hbfe4397f5b2a4380, 64'h3fe8cc6a75184655,
	64'h3fb9dfb6eb24a85c, 64'h3fefd60d2da75c9e,
	64'hbfefd60d2da75c9e, 64'h3fb9dfb6eb24a85c,
	64'h3fef677556883cee, 64'h3fc8961727c41804,
	64'hbfc8961727c41804, 64'h3fef677556883cee,
	64'h3fe1dc1b64dc4872, 64'h3fea8d676e545ad2,
	64'hbfea8d676e545ad2, 64'h3fe1dc1b64dc4872,
	64'h3feaa9547a2cb98e, 64'h3fe1b250171373bf,
	64'hbfe1b250171373bf, 64'h3feaa9547a2cb98e,
	64'h3fc95b49e9b62afa, 64'h3fef5da6ed43685d,
	64'hbfef5da6ed43685d, 64'h3fc95b49e9b62afa,
	64'h3fed9a00dd8b3d46, 64'h3fd84f6aaaf3903f,
	64'hbfd84f6aaaf3903f, 64'h3fed9a00dd8b3d46,
	64'h3fd8ac4b86d5ed44, 64'h3fed86c48445a44f,
	64'hbfed86c48445a44f, 64'h3fd8ac4b86d5ed44,
	64'h3fe6b25ced2fe29c, 64'h3fe68ed1eaa19c71,
	64'hbfe68ed1eaa19c71, 64'h3fe6b25ced2fe29c,
	64'h3f6921f8becca4ba, 64'h3feffff621621d02,
	64'hbfeffff621621d02, 64'h3f6921f8becca4ba
};

//---------------------------------------------------------------------
//   REG & WIRE DECLARATION
//---------------------------------------------------------------------
reg [FLOAT_PRECISION-1:0] f_re [0:n-1], f_im[0:n-1];
reg [FLOAT_PRECISION-1:0] s_index [0:n-1];
reg [FLOAT_PRECISION-1:0] golden_fo_re [0:n-1], golden_fo_im [0:n-1];
reg [FLOAT_PRECISION-1:0] your_fo_re [0:n-1], your_fo_im [0:n-1];

//---------------------------------------------------------------------
//   Clock
//---------------------------------------------------------------------
real CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;

//---------------------------------------------------------------------
//  Simulation
//---------------------------------------------------------------------
initial begin
	file_in = $fopen(INPUT_PATH, "r");
	file_idx = $fopen(INDEX_PATH, "r");
	file_out = $fopen(OUTPUT_PATH, "r");
	file_num = $fopen(PATNUM_PATH, "r");
	fscanf_int = $fscanf(file_num, "%d", PAT_NUM);	

	reset_task;
	total_latency = 0;
	repeat(4) @(negedge clk);
	for (i_pat = 0; i_pat < PAT_NUM; i_pat = i_pat + 1)begin
		read_pattern;
		i_in_deg = 0;
		i_out_deg = 0;
		pattern_latency = 0;
		while (i_in_deg < n) begin
			input_task;
			if (i_in_deg != n)
				input_delay;
		end		
		in_valid = 'b0;
		fi_re = 'bx;
		fi_im = 'bx;
		while (i_out_deg < n) begin
			@(negedge clk);		
			in_valid = 'b0;
			wait_out_task;
			pattern_latency = pattern_latency + out_latency;			
			total_latency = total_latency + out_latency;
		end
		$display("PASS PATTERN NO.%4d, %4d CYCLES", i_pat+1, pattern_latency);
		repeat($urandom_range(2, 4)) @(negedge clk);
	end
	YOU_PASS_task;
end

always @(negedge clk) begin
	check_ans_task;
	twiddle_factor;
end

//---------------------------------------------------------------------
//   Task
//---------------------------------------------------------------------
task reset_task; begin 
    rst_n = 'b1;
    in_valid = 'b0;
    fi_re = 'bx;
    fi_im = 'bx;
    s_re_1 = 'bx; s_im_1 = 'bx;
    s_re_2 = 'bx; s_im_2 = 'bx;
    s_re_3 = 'bx; s_im_3 = 'bx;
    s_re_4 = 'bx; s_im_4 = 'bx;
    s_re_5 = 'bx; s_im_5 = 'bx;
    s_re_6 = 'bx; s_im_6 = 'bx;
    s_re_7 = 'bx; s_im_7 = 'bx;
    s_re_8 = 'bx; s_im_8 = 'bx;
	
    force clk = 0;
    #CYCLE; rst_n = 0; 
    #CYCLE; rst_n = 1;
    if(out_valid !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'out_valid' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_1 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_1' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_2 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_2' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_3 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_3' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_4 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_4' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_5 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_5' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_6 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_6' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_7 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_7' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(tw_idx_8 !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'tw_idx_8' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(fo_re !== 'b0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'fo_re' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
    if(fo_im !== 0) begin 
        $display("************************************************************");  
        $display("                          FAIL!                             ");    
        $display("  'fo_im' should be 0 after initial RESET  at %8t   	  ",$time);
        $display("************************************************************");
        repeat(2) #CYCLE;
        $finish;
    end
	#CYCLE; release clk;
end endtask


task read_pattern; begin
	for (i_in_deg = 0; i_in_deg < n; i_in_deg = i_in_deg + 1) 
		fscanf_int = $fscanf(file_in, "%h", f_re[i_in_deg]);
	for (i_in_deg = 0; i_in_deg < n; i_in_deg = i_in_deg + 1) 
		fscanf_int = $fscanf(file_in, "%h", f_im[i_in_deg]);
	for (i_in_deg = 0; i_in_deg < n; i_in_deg = i_in_deg + 1) 
		fscanf_int = $fscanf(file_out, "%h", golden_fo_re[i_in_deg]);
	for (i_in_deg = 0; i_in_deg < n; i_in_deg = i_in_deg + 1) 
		fscanf_int = $fscanf(file_out, "%h", golden_fo_im[i_in_deg]);
	for (i_in_deg = 0; i_in_deg < n; i_in_deg = i_in_deg + 1) 
		fscanf_int = $fscanf(file_idx, "%d", s_index[i_in_deg]);
end endtask

task input_task; begin
	in_valid = 'b1;
	fi_re = f_re[i_in_deg];
	fi_im = f_im[i_in_deg];
	// $display("\tIN  DEGREE %3d\tRe = %f, Im = %f", i_in_deg, $bitstoreal(fi_re), $bitstoreal(fi_im));
	i_in_deg = i_in_deg + 1;
	@(negedge clk);		
end endtask

task twiddle_factor; begin
	s_re_1 = fpr_gm_tab[(tw_idx_1 << 1) + 0];
	s_im_1 = fpr_gm_tab[(tw_idx_1 << 1) + 1];
	s_re_2 = fpr_gm_tab[(tw_idx_2 << 1) + 0];
	s_im_2 = fpr_gm_tab[(tw_idx_2 << 1) + 1];
	s_re_3 = fpr_gm_tab[(tw_idx_3 << 1) + 0];
	s_im_3 = fpr_gm_tab[(tw_idx_3 << 1) + 1];
	s_re_4 = fpr_gm_tab[(tw_idx_4 << 1) + 0];
	s_im_4 = fpr_gm_tab[(tw_idx_4 << 1) + 1];
	s_re_5 = fpr_gm_tab[(tw_idx_5 << 1) + 0];
	s_im_5 = fpr_gm_tab[(tw_idx_5 << 1) + 1];
	s_re_6 = fpr_gm_tab[(tw_idx_6 << 1) + 0];
	s_im_6 = fpr_gm_tab[(tw_idx_6 << 1) + 1];
	s_re_7 = fpr_gm_tab[(tw_idx_7 << 1) + 0];
	s_im_7 = fpr_gm_tab[(tw_idx_7 << 1) + 1];
	s_re_8 = fpr_gm_tab[(tw_idx_8 << 1) + 0];
	s_im_8 = fpr_gm_tab[(tw_idx_8 << 1) + 1];
	// $display("s1: Re = %f, Im = %f", $bitstoreal(s_re_1), $bitstoreal(s_im_1));
	// $display("s2 (%3d): Re = %f, Im = %f", tw_idx_2, $bitstoreal(s_re_2), $bitstoreal(s_im_2));
end endtask

task input_delay; begin
	integer DELAY_NUM;
	DELAY_NUM = $urandom_range(1, 4);
	// DELAY_NUM = 0;
	for (i_delay = 0; i_delay < DELAY_NUM; i_delay=i_delay+1) begin
		in_valid = 'b0;
		fi_re = 'bx;
		fi_im = 'bx;
		@(negedge clk);
end
end endtask

task wait_out_task; begin
	out_latency = 1;
	while(out_valid !== 1 && i_out_deg < n) begin
		if(out_latency === MAX_OUT_LATENCY + 1) begin
            $display("***********************************************************");    
            $display("                          FAIL!                          	 ");
			$display("         The execution latency are over %d cycles        	 ", MAX_OUT_LATENCY);
		    $display("***********************************************************"); 
			repeat(2) @(negedge clk);
			$finish;
		end
		out_latency = out_latency + 1;
		@(negedge clk);
	end
end endtask

task check_out_valid_task; begin
	if(out_valid !== 0) begin
		$display("***********************************************************");     
        $display("*                          FAIL!                          *");
		$display("*  out_valid should not be raised when in_valid is high.  *");
		$display("***********************************************************");
		repeat(2) @(negedge clk);
		$finish;
	end
end endtask

task check_ans_task; begin
	if(out_valid == 1) begin
		// $display("\tOUT DEGREE %3d\tRe = %f, Im = %f", i_out_deg, $bitstoreal(golden_fo_re[i_out_deg]), $bitstoreal(golden_fo_im[i_out_deg]));
		if(fo_re !== golden_fo_re[i_out_deg] || fo_im !== golden_fo_im[i_out_deg])begin
            $display("***********************************************************");     
            $display("                          FAIL!                          	 ");  
            $display("                  Degree #%3d (%8t)                   	 ", i_out_deg, $time);
            $display("                      Golden answer                      	 ");
            $display("              Re = %f, Im = %f                    	     ", $bitstoreal(golden_fo_re[i_out_deg]), $bitstoreal(golden_fo_im[i_out_deg]));
            $display("                       Your answer                       	 ");
            $display("              Re = %f, Im = %f                    	     ", $bitstoreal(fo_re), $bitstoreal(fo_im));
            $display("***********************************************************");    
                repeat(2) @(negedge clk);
                $finish;
		end
		i_out_deg = i_out_deg + 1;
	end
end endtask

task YOU_PASS_task; begin
    $display ("--------------------------------------------------------------------");
    $display ("                         Congratulations!                           ");
    $display ("                  You have passed all patterns!                     ");
    $display ("                  Your execution cycles = %5d cycles                ", total_latency);
	$display ("                  Your clock period = %.1f ns                       ", CYCLE);
    $display ("                  Total Latency = %.1f ns                           ", total_latency*CYCLE);
    $display ("--------------------------------------------------------------------");     
    repeat(2)@(negedge clk);
    $finish;
end endtask

endmodule