//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM, INC.
//Copyright (c) 2002-2009 ARM, Inc.
//The confidential and proprietary information contained in this file
//may only be used by a person authorised under and to the extent
//permitted by a subsisting licensing agreement from ARM Limited.
//
//(C) COPYRIGHT 2004-2009 ARM Limited.
//ALL RIGHTS RESERVED
//
//This entire notice must be reproduced on all copies of this file
//and copies of this file may only be made by a person if such person
//is permitted to do so under the terms of a subsisting license
//agreement from ARM Limited.
//

`ifdef ARM_UD_MODEL

`ifdef ARM_UD_DP
`else
`define ARM_UD_DP #0.001
`endif
`ifdef ARM_UD_CP
`else
`define ARM_UD_CP
`endif
`ifdef ARM_UD_SEQ
`else
`define ARM_UD_SEQ #0.01
`endif

`timescale 1ns/1ps

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X0P5M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // A2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X1M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // A2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X2M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // A2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X3M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // A2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X0P5M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // A2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X1M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // A2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X2M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // A2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X3M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // A2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X4M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // A2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or `ARM_UD_DP I5 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1P4M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or `ARM_UD_DP I5 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X2M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or `ARM_UD_DP I5 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1P4M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X2M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1P4M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X2M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1P4M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X2M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X11M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X8M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X6M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X8M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4_X8M_A9TH
`endcelldefine
module ANTENNA1_A9TH (A);
input A;

endmodule // ANTENNA1_A9TH

`timescale 1ns/1ps
`celldefine
module AO1B2_X0P5M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X0P7M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1P4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X2M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X3M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X6M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // AO1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand `ARM_UD_DP I3(Y, outB, C0);


endmodule // AO21A1AI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or `ARM_UD_DP I2(Y, outB, outA);
endmodule // AO21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or `ARM_UD_DP I1(Y, B0, outA);
endmodule // AO21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or `ARM_UD_DP I2(Y, outA, outB);
endmodule // AO22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor `ARM_UD_DP I3 (Y,outA,outB);
endmodule // AOI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P5M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P7M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1P4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X2M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X3M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P5M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P7M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1P4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X2M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X3M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P5M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P7M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1P4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X2M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X3M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X6M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X8M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor `ARM_UD_DP I4 (Y,outA,outB);
endmodule // AOI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P5M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P7M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1P4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X2M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X3M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X6M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X8M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor `ARM_UD_DP I2(Y, B0, outA);
endmodule // AOI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P5M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P7M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1P4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X2M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X3M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X6M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P5M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P7M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1P4M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X2M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X3M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X4M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X6M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X11M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X16M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X2M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X3M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X4M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X6M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X8M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENC_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X0P7M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  `ARM_UD_DP I1 (PPN, nPP);

endmodule // BMXIT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  `ARM_UD_DP I1 (PPN, nPP);

endmodule // BMXIT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1P4M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  `ARM_UD_DP I1 (PPN, nPP);

endmodule // BMXIT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X2M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  `ARM_UD_DP I1 (PPN, nPP);

endmodule // BMXIT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X0P7M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx `ARM_UD_DP I0 (PP, X2, AN, SN, D1, D0);

endmodule // BMXT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx `ARM_UD_DP I0 (PP, X2, AN, SN, D1, D0);

endmodule // BMXT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1P4M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx `ARM_UD_DP I0 (PP, X2, AN, SN, D1, D0);

endmodule // BMXT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X2M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx `ARM_UD_DP I0 (PP, X2, AN, SN, D1, D0);

endmodule // BMXT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P7M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P8M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X11M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X13M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X16M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P2M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P4M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P7M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X4M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X6M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X7P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X9M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFH_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X11M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X16M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1P4M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X2M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X3M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X4M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X6M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X8M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // BUFZ_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUF_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGENCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1P4M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGENCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X2M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGENCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENCON_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1P4M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENCON_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X2M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENCON_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1P4M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENI_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X2M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I4 (CON, cout);
endmodule // CGENI_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGEN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1P4M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGEN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X2M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or `ARM_UD_DP I4 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // CGEN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  `ARM_UD_DP  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor `ARM_UD_DP  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  `ARM_UD_DP  I11 (CO, t5, t6, t7);

endmodule // CMPR42_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1P4M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  `ARM_UD_DP  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor `ARM_UD_DP  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  `ARM_UD_DP  I11 (CO, t5, t6, t7);

endmodule // CMPR42_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X2M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  `ARM_UD_DP  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor `ARM_UD_DP  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  `ARM_UD_DP  I11 (CO, t5, t6, t7);

endmodule // CMPR42_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFNQ_X1M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X2M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X3M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X1M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X2M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X3M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFNSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X0P5M_A9TH (QN, CK, D);
output QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X1M_A9TH (QN, CK, D);
output QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X2M_A9TH (QN, CK, D);
output QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X3M_A9TH (QN, CK, D);
output QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X0P5M_A9TH (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X1M_A9TH (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X2M_A9TH (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X3M_A9TH (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X4M_A9TH (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X0P5M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRPQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X1M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRPQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X2M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRPQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X3M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRPQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X0P5M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X1M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X2M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X3M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X4M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
supply1 xSN;

  not   XX0 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X0P5M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X1M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X2M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X3M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X0P5M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X1M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X2M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X3M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X4M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff I0 (n0, D, CK, xRN, SN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X0P5M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X1M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X2M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X3M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X4M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  udp_dff I0 (n0, D, CK, xRN, xSN, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY2_X0P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // DLY2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X1M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // DLY2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X0P5M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // DLY4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X1M_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // DLY4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S2_X1B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // DLYCLK8S2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S4_X1B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // DLYCLK8S4_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S6_X1B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // DLYCLK8S6_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S8_X1B_A9TH ( Y, A );
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // DLYCLK8S8_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ENDCAPTIE3_A9TH;

endmodule // ENDCAPTIE3_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ESDFFQN_X0P5M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   not       `ARM_UD_SEQ I1 (QN, n0);
endmodule // ESDFFQN_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X1M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   not       `ARM_UD_SEQ I1 (QN, n0);
endmodule // ESDFFQN_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X2M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   not       `ARM_UD_SEQ I1 (QN, n0);
endmodule // ESDFFQN_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X3M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   not       `ARM_UD_SEQ I1 (QN, n0);
endmodule // ESDFFQN_X3M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X0P5M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // ESDFFQ_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X1M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // ESDFFQ_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X2M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // ESDFFQ_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X3M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // ESDFFQ_X3M_A9TH
`endcelldefine


module FILL128_A9TH;

endmodule // FILL128_A9TH

module FILL16_A9TH;

endmodule // FILL16_A9TH

module FILL1_A9TH;

endmodule // FILL1_A9TH

module FILL2_A9TH;

endmodule // FILL2_A9TH

module FILL32_A9TH;

endmodule // FILL32_A9TH

module FILL4_A9TH;

endmodule // FILL4_A9TH

module FILL64_A9TH;

endmodule // FILL64_A9TH

module FILL8_A9TH;

endmodule // FILL8_A9TH

module FILLCAP128_A9TH;

endmodule // FILLCAP128_A9TH

module FILLCAP16_A9TH;

endmodule // FILLCAP16_A9TH

module FILLCAP32_A9TH;

endmodule // FILLCAP32_A9TH

module FILLCAP4_A9TH;

endmodule // FILLCAP4_A9TH

module FILLCAP64_A9TH;

endmodule // FILLCAP64_A9TH

module FILLCAP8_A9TH;

endmodule // FILLCAP8_A9TH

module FILLSGCAP128_A9TH;

endmodule // FILLSGCAP128_A9TH

module FILLSGCAP16_A9TH;

endmodule // FILLSGCAP16_A9TH

module FILLSGCAP32_A9TH;

endmodule // FILLSGCAP32_A9TH

module FILLSGCAP4_A9TH;

endmodule // FILLSGCAP4_A9TH

module FILLSGCAP64_A9TH;

endmodule // FILLSGCAP64_A9TH

module FILLSGCAP8_A9TH;

endmodule // FILLSGCAP8_A9TH

module FILLTIE128_A9TH;

endmodule // FILLTIE128_A9TH

module FILLTIE16_A9TH;

endmodule // FILLTIE16_A9TH

module FILLTIE32_A9TH;

endmodule // FILLTIE32_A9TH

module FILLTIE3_A9TH;

endmodule // FILLTIE3_A9TH

module FILLTIE4_A9TH;

endmodule // FILLTIE4_A9TH

module FILLTIE64_A9TH;

endmodule // FILLTIE64_A9TH

module FILLTIE8_A9TH;

endmodule // FILLTIE8_A9TH

`timescale 1ns/1ps
`celldefine
module FRICG_X0P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P6B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P7B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P8B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X11B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X13B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X16B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P2B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P4B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P7B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X4B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X6B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X7P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X9B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf `ARM_UD_DP I0(ECK, CK);

endmodule // FRICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9B_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9M_A9TH ( Y, A );
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INV_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X0P5M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X1M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X2M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X3M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X4M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X0P5M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X1M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X2M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X3M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X0P5M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X1M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X2M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X3M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X4M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X0P5M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, GN, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X1M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, GN, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X2M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, GN, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X3M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, GN, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X0P5M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X1M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X2M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X3M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, GN, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
buf      I3 (clk, GN);
endmodule // LATNSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X0P5M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, GN, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X1M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, GN, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X2M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, GN, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X3M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, GN, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X4M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, GN, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // LATNSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X0P5M_A9TH (QN, D, G);
output  QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X1M_A9TH (QN, D, G);
output  QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X2M_A9TH (QN, D, G);
output  QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X3M_A9TH (QN, D, G);
output  QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X4M_A9TH (QN, D, G);
output  QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X0P5M_A9TH (Q, D, G);
output  Q;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X1M_A9TH (Q, D, G);
output  Q;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X2M_A9TH (Q, D, G);
output  Q;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X3M_A9TH (Q, D, G);
output  Q;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X0P5M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X1M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X2M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X3M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X4M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X0P5M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, clk, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X1M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, clk, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X2M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, clk, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X3M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat I0 (n0, D, clk, RN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X0P5M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X1M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X2M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X3M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not  I3(clk,G);
endmodule // LATSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X0P5M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, clk, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X1M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, clk, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X2M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, clk, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X3M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, clk, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X4M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat I0 (n0, D, clk, xRN, SN, 1'b1);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // LATSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X0P5M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // M2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X1M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // M2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X2M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // M2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X3M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  not     `ARM_UD_SEQ I3 (QN, n0);
endmodule // M2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X0P5M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // M2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X1M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // M2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X2M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // M2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X3M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // M2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X4M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I2 (n1, nm, SI, SE);
  buf     `ARM_UD_SEQ I3 (Q, n0);
endmodule // M2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module MX2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X8B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXGL2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P5M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P7M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1P4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X2M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X3M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P5M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P7M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1P4M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X2M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X3M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXIT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MXT2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P5M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P7M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1P4M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X2M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X3M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MXT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P5M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P7M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1P4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X2M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X3M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X6M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X8M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P5M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P7M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1P4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X2M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X3M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X6M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X8M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand `ARM_UD_DP (Y, A, Bx);
endmodule // NAND2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8A_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P5M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P7M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1P4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X2M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X3M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X6M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X8M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NAND3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P5M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P7M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1P4M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X2M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X3M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X4M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X6M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P5M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P7M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1P4M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X2M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X3M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X4M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X6M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand `ARM_UD_DP (Y, A, B, Cx);
endmodule // NAND3XXB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P5M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P7M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1P4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X2M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X3M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X6M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P5M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P7M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1P4M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X2M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X3M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X4M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P5M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P7M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1P4M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X2M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X3M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X4M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand `ARM_UD_DP (Y, A, B, C, Dx);
endmodule // NAND4XXXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P5M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P7M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1P4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X2M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X3M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X6M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X8M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P5M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P7M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1P4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X2M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X3M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X6M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X8M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor `ARM_UD_DP (Y, A, Bx);
endmodule // NOR2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8A_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P5M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P7M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1P4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X2M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X3M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X6M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X8M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C);
endmodule // NOR3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P5M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P7M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1P4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X2M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X3M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P5M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P7M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1P4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X2M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X3M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X6M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X8M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor `ARM_UD_DP I2 (Y, A0N, outB);
endmodule // OA1B2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OA211_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor `ARM_UD_DP I3(Y, outB, C0);

endmodule // OA21A1OI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and `ARM_UD_DP I2(Y, outB, outA);
endmodule // OA21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and `ARM_UD_DP I1(Y, B0, outA);
endmodule // OA21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and `ARM_UD_DP I2(Y, outA, outB);
endmodule // OA22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand `ARM_UD_DP I2 (Y, outA, outB);
endmodule // OAI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P5M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P7M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1P4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X2M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X3M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P5M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P7M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1P4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X2M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X3M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P5M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P7M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1P4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X2M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X3M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X6M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X8M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand `ARM_UD_DP I4 (Y, outA, outB);
endmodule // OAI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P5M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P7M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1P4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X2M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X3M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X6M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X8M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand `ARM_UD_DP I2 (Y, B0, outA);
endmodule // OAI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P5M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P7M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1P4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X2M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X3M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X6M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X8M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X6M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X8M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P5M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P7M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1P4M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X2M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X3M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X4M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X6M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or `ARM_UD_DP (Y, A, B, C, D, E, F);
endmodule // OR6_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P6B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P7B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P8B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X11B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X13B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X16B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P2B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P4B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P7B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X4B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X6B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X7P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X9B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // POSTICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P6B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P7B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P8B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X11B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X13B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X16B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P2B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P4B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P7B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X4B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X6B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X7P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X9B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // PREICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  1'b1);
   bufif1     `ARM_UD_SEQ I1 (RBL, n0, RWL);




endmodule // RF1R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1P4M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  1'b1);
   bufif1     `ARM_UD_SEQ I1 (RBL, n0, RWL);




endmodule // RF1R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X2M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  1'b1);
   bufif1     `ARM_UD_SEQ I1 (RBL, n0, RWL);




endmodule // RF1R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1  `ARM_UD_SEQ  I5(RBL, n1, RWL);




endmodule // RF1R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1P4M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1  `ARM_UD_SEQ  I5(RBL, n1, RWL);




endmodule // RF1R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X2M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1  `ARM_UD_SEQ  I5(RBL, n1, RWL);




endmodule // RF1R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  1'b1);
   bufif1     `ARM_UD_SEQ I4 (RBL1, n0, n2);
   bufif1     `ARM_UD_SEQ I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);




endmodule // RF2R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1P4M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  1'b1);
   bufif1     `ARM_UD_SEQ I4 (RBL1, n0, n2);
   bufif1     `ARM_UD_SEQ I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);




endmodule // RF2R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X2M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  1'b1);
   bufif1     `ARM_UD_SEQ I4 (RBL1, n0, n2);
   bufif1     `ARM_UD_SEQ I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);




endmodule // RF2R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1 `ARM_UD_SEQ I5 (RBL1, n1, RWL1);
   bufif1 `ARM_UD_SEQ I6 (RBL2, n1, RWL2);




endmodule // RF2R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1P4M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1 `ARM_UD_SEQ I5 (RBL1, n1, RWL1);
   bufif1 `ARM_UD_SEQ I6 (RBL2, n1, RWL2);




endmodule // RF2R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X2M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 `ARM_UD_SEQ I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, 1'b1);
   not I4 (n1, n0);
   bufif1 `ARM_UD_SEQ I5 (RBL1, n1, RWL1);
   bufif1 `ARM_UD_SEQ I6 (RBL2, n1, RWL2);




endmodule // RF2R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFNQ_X1M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X2M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X3M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X1M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X2M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X3M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X1M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X2M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X3M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X1M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X2M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X3M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFNSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X0P5M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X1M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X2M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X3M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X0P5M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X1M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X2M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X3M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X4M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X0P5M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRPQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X1M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRPQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X2M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRPQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X3M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRPQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X0P5M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X1M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X2M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X3M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X4M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X0P5M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X1M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X2M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X3M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X0P5M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X1M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X2M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X3M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X4M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff I0 (n0, n1, CK, xRN, SN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X0P5M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X1M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X2M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X3M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X4M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X1M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFYQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X2M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFYQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X3M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFYQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X4M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff I0 (n0, n1, CK, xRN, xSN, 1'b1);
  udp_mux I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFYQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module TIEHI_X1M_A9TH (Y);
output Y;

  buf I0(Y, 1'b1);

endmodule // TIEHI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO_X1M_A9TH (Y);
output Y;

  buf I0(Y, 1'b0);

endmodule // TIELO_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3_X4M_A9TH
`endcelldefine
`else

`define ARM_PROP_DELAY 1.0
`define ARM_PERIOD 1.0
`define ARM_WIDTH 1.0
`define ARM_SETUP_TIME 1.0
`define ARM_HOLD_TIME 0.5
`define ARM_RECOVERY_TIME 1.0
`define ARM_REMOVAL_TIME 0.5

`timescale 1ns/1ps

`ifdef POWER_PINS
`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X0P5M_A9TH (QN,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X1M_A9TH (QN,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X2M_A9TH (QN,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X3M_A9TH (QN,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X0P5M_A9TH (Q,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X1M_A9TH (Q,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X2M_A9TH (Q,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X3M_A9TH (Q,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X4M_A9TH (Q,VDD, VSS, A, B, CK, SE, SI);
inout VDD, VSS;
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1M_A9TH ( CO, SUM,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, B, ci);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1P4M_A9TH ( CO, SUM,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, B, ci);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X2M_A9TH ( CO, SUM,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, B, ci);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1M_A9TH ( CO, SUM,VDD, VSS, A, B, CI);
inout VDD, VSS;
output SUM, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1P4M_A9TH ( CO, SUM,VDD, VSS, A, B, CI);
inout VDD, VSS;
output SUM, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X2M_A9TH ( CO, SUM,VDD, VSS, A, B, CI);
inout VDD, VSS;
output SUM, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1M_A9TH ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1P4M_A9TH ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X2M_A9TH ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1M_A9TH ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1P4M_A9TH ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X2M_A9TH ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X11M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X6M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X8M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X2M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X3M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X6M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X8M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X8M_A9TH
`endcelldefine
module ANTENNA1_A9TH (A,VDD, VSS);
inout VDD, VSS;
input A;


specify

endspecify
endmodule // ANTENNA1_A9TH
`timescale 1ns/1ps
`celldefine
module AO1B2_X0P5M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X0P7M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1P4M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X2M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X3M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X4M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X6M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X2M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X3M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X6M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X8M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X2M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X3M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X6M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X8M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X8M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X8M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P5M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P7M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1P4M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X2M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X3M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X4M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X6M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X8M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P5M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P7M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1P4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X2M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X3M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X6M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P5M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P7M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1P4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X2M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X3M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X6M_A9TH (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X11M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X16M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X2M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X3M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X4M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X6M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X8M_A9TH (AN, SN, X2,VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign SN = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign AN = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X0P7M_A9TH (PPN,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN_temp, nPP);
  assign PPN = ((VDD === 1'b1) && (VSS === 1'b0))? PPN_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1M_A9TH (PPN,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN_temp, nPP);
  assign PPN = ((VDD === 1'b1) && (VSS === 1'b0))? PPN_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1P4M_A9TH (PPN,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN_temp, nPP);
  assign PPN = ((VDD === 1'b1) && (VSS === 1'b0))? PPN_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X2M_A9TH (PPN,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN_temp, nPP);
  assign PPN = ((VDD === 1'b1) && (VSS === 1'b0))? PPN_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X0P7M_A9TH (PP,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (z_temp, X2, AN, SN, D1, D0);
  assign PP = ((VDD === 1'b1) && (VSS === 1'b0))? z_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1M_A9TH (PP,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (z_temp, X2, AN, SN, D1, D0);
  assign PP = ((VDD === 1'b1) && (VSS === 1'b0))? z_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1P4M_A9TH (PP,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (z_temp, X2, AN, SN, D1, D0);
  assign PP = ((VDD === 1'b1) && (VSS === 1'b0))? z_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X2M_A9TH (PP,VDD, VSS, AN, D0, D1, SN, X2);
inout VDD, VSS;
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (z_temp, X2, AN, SN, D1, D0);
  assign PP = ((VDD === 1'b1) && (VSS === 1'b0))? z_temp : 1'bx;



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P8M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X11M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X13M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X16M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X6M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X7P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X9M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X11M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X16M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1P4M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X2M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X3M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X4M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X6M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X8M_A9TH ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1M_A9TH ( CO,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1P4M_A9TH ( CO,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X2M_A9TH ( CO,VDD, VSS, A, B, CIN);
inout VDD, VSS;
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1P4M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X2M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1P4M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X2M_A9TH ( CON,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1M_A9TH ( CO,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1P4M_A9TH ( CO,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X2M_A9TH ( CO,VDD, VSS, A, B, CI);
inout VDD, VSS;
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1M_A9TH (CO, ICO, SUM,VDD, VSS, A, B, C, D, ICI);
inout VDD, VSS;
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (co_temp, t2, t3, t4);
  assign ICO = ((VDD === 1'b1) && (VSS === 1'b0))? co_temp : 1'bx;
  xor I6 (ss, IS, D);
  xor  I7 (sum_temp, ss, ICI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (c_temp, t5, t6, t7);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? c_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1P4M_A9TH (CO, ICO, SUM,VDD, VSS, A, B, C, D, ICI);
inout VDD, VSS;
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (co_temp, t2, t3, t4);
  assign ICO = ((VDD === 1'b1) && (VSS === 1'b0))? co_temp : 1'bx;
  xor I6 (ss, IS, D);
  xor  I7 (sum_temp, ss, ICI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (c_temp, t5, t6, t7);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? c_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X2M_A9TH (CO, ICO, SUM,VDD, VSS, A, B, C, D, ICI);
inout VDD, VSS;
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (co_temp, t2, t3, t4);
  assign ICO = ((VDD === 1'b1) && (VSS === 1'b0))? co_temp : 1'bx;
  xor I6 (ss, IS, D);
  xor  I7 (sum_temp, ss, ICI);
  assign SUM = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (c_temp, t5, t6, t7);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? c_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFNQ_X1M_A9TH (Q,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X2M_A9TH (Q,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X3M_A9TH (Q,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X1M_A9TH (Q,VDD, VSS, CKN, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X2M_A9TH (Q,VDD, VSS, CKN, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X3M_A9TH (Q,VDD, VSS, CKN, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X0P5M_A9TH (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X1M_A9TH (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X2M_A9TH (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X3M_A9TH (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X0P5M_A9TH (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X1M_A9TH (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X2M_A9TH (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X3M_A9TH (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X4M_A9TH (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, R);
inout VDD, VSS;
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X1M_A9TH (QN,VDD, VSS, CK, D, R);
inout VDD, VSS;
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X2M_A9TH (QN,VDD, VSS, CK, D, R);
inout VDD, VSS;
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X3M_A9TH (QN,VDD, VSS, CK, D, R);
inout VDD, VSS;
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, R);
inout VDD, VSS;
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X1M_A9TH (Q,VDD, VSS, CK, D, R);
inout VDD, VSS;
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X2M_A9TH (Q,VDD, VSS, CK, D, R);
inout VDD, VSS;
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X3M_A9TH (Q,VDD, VSS, CK, D, R);
inout VDD, VSS;
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X4M_A9TH (Q,VDD, VSS, CK, D, R);
inout VDD, VSS;
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X1M_A9TH (QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X2M_A9TH (QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X3M_A9TH (QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X1M_A9TH (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X2M_A9TH (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X3M_A9TH (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X4M_A9TH (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X1M_A9TH (Q,VDD, VSS, CK, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X2M_A9TH (Q,VDD, VSS, CK, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X3M_A9TH (Q,VDD, VSS, CK, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X4M_A9TH (Q,VDD, VSS, CK, D, R, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY2_X0P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X1M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X0P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X1M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S2_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S4_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S4_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S6_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S6_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S8_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S8_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ENDCAPTIE3_A9TH (VDD, VSS);
inout VDD, VSS;

endmodule //ENDCAPTIE3_A9TH

`endcelldefine
`timescale 1ns/1ps
`celldefine
module ESDFFQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   not       I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X1M_A9TH (QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   not       I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X2M_A9TH (QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   not       I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X3M_A9TH (QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   not       I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X3M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X1M_A9TH (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X2M_A9TH (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X3M_A9TH (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X3M_A9TH
`endcelldefine


module FILL128_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL128_A9TH

module FILL16_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL16_A9TH

module FILL1_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL1_A9TH

module FILL2_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL2_A9TH

module FILL32_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL32_A9TH

module FILL4_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL4_A9TH

module FILL64_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL64_A9TH

module FILL8_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILL8_A9TH

module FILLCAP128_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP128_A9TH
module FILLCAP16_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP16_A9TH
module FILLCAP32_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP32_A9TH
module FILLCAP4_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP4_A9TH
module FILLCAP64_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP64_A9TH
module FILLCAP8_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP8_A9TH
module FILLSGCAP128_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP128_A9TH
module FILLSGCAP16_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP16_A9TH
module FILLSGCAP32_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP32_A9TH
module FILLSGCAP4_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP4_A9TH
module FILLSGCAP64_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP64_A9TH
module FILLSGCAP8_A9TH (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLSGCAP8_A9TH
module FILLTIE128_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE128_A9TH

module FILLTIE16_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE16_A9TH

module FILLTIE32_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE32_A9TH

module FILLTIE3_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE3_A9TH

module FILLTIE4_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE4_A9TH

module FILLTIE64_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE64_A9TH

module FILLTIE8_A9TH (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE8_A9TH

`timescale 1ns/1ps
`celldefine
module FRICG_X0P5B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P6B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P7B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P8B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X11B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X13B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X16B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P2B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P4B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P7B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2P5B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3P5B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X4B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X5B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X6B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X7P5B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X9B_A9TH ( ECK,VDD, VSS, CK );
inout VDD, VSS;
output ECK;
input CK;

  buf I0(out_temp, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9B_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9M_A9TH ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X0P5M_A9TH (QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X1M_A9TH (QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X2M_A9TH (QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X3M_A9TH (QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X4M_A9TH (QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X0P5M_A9TH (Q,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X1M_A9TH (Q,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X2M_A9TH (Q,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X3M_A9TH (Q,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X0P5M_A9TH (QN,VDD, VSS, D, GN, R);
inout VDD, VSS;
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X1M_A9TH (QN,VDD, VSS, D, GN, R);
inout VDD, VSS;
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X2M_A9TH (QN,VDD, VSS, D, GN, R);
inout VDD, VSS;
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X3M_A9TH (QN,VDD, VSS, D, GN, R);
inout VDD, VSS;
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X4M_A9TH (QN,VDD, VSS, D, GN, R);
inout VDD, VSS;
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X0P5M_A9TH (Q,VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X1M_A9TH (Q,VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X2M_A9TH (Q,VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X3M_A9TH (Q,VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X0P5M_A9TH (Q,VDD, VSS, D, GN, S);
inout VDD, VSS;
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X1M_A9TH (Q,VDD, VSS, D, GN, S);
inout VDD, VSS;
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X2M_A9TH (Q,VDD, VSS, D, GN, S);
inout VDD, VSS;
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X3M_A9TH (Q,VDD, VSS, D, GN, S);
inout VDD, VSS;
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X0P5M_A9TH (QN,VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X1M_A9TH (QN,VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X2M_A9TH (QN,VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X3M_A9TH (QN,VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X4M_A9TH (QN,VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X0P5M_A9TH (QN,VDD, VSS, D, G);
inout VDD, VSS;
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X1M_A9TH (QN,VDD, VSS, D, G);
inout VDD, VSS;
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X2M_A9TH (QN,VDD, VSS, D, G);
inout VDD, VSS;
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X3M_A9TH (QN,VDD, VSS, D, G);
inout VDD, VSS;
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X4M_A9TH (QN,VDD, VSS, D, G);
inout VDD, VSS;
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X0P5M_A9TH (Q,VDD, VSS, D, G);
inout VDD, VSS;
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X1M_A9TH (Q,VDD, VSS, D, G);
inout VDD, VSS;
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X2M_A9TH (Q,VDD, VSS, D, G);
inout VDD, VSS;
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X3M_A9TH (Q,VDD, VSS, D, G);
inout VDD, VSS;
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X0P5M_A9TH (QN,VDD, VSS, D, G, R);
inout VDD, VSS;
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X1M_A9TH (QN,VDD, VSS, D, G, R);
inout VDD, VSS;
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X2M_A9TH (QN,VDD, VSS, D, G, R);
inout VDD, VSS;
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X3M_A9TH (QN,VDD, VSS, D, G, R);
inout VDD, VSS;
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X4M_A9TH (QN,VDD, VSS, D, G, R);
inout VDD, VSS;
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X0P5M_A9TH (Q,VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X1M_A9TH (Q,VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X2M_A9TH (Q,VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X3M_A9TH (Q,VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X0P5M_A9TH (Q,VDD, VSS, D, G, S);
inout VDD, VSS;
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X1M_A9TH (Q,VDD, VSS, D, G, S);
inout VDD, VSS;
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X2M_A9TH (Q,VDD, VSS, D, G, S);
inout VDD, VSS;
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X3M_A9TH (Q,VDD, VSS, D, G, S);
inout VDD, VSS;
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X0P5M_A9TH (QN,VDD, VSS, D, G, SN);
inout VDD, VSS;
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X1M_A9TH (QN,VDD, VSS, D, G, SN);
inout VDD, VSS;
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X2M_A9TH (QN,VDD, VSS, D, G, SN);
inout VDD, VSS;
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X3M_A9TH (QN,VDD, VSS, D, G, SN);
inout VDD, VSS;
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X4M_A9TH (QN,VDD, VSS, D, G, SN);
inout VDD, VSS;
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X0P5M_A9TH (QN,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X1M_A9TH (QN,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X2M_A9TH (QN,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X3M_A9TH (QN,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X0P5M_A9TH (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X1M_A9TH (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X2M_A9TH (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X3M_A9TH (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X4M_A9TH (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff_PWR  I1 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module MX2_X0P5B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X0P7B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1P4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X2B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X3B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X6B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X8B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P5B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P7B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1P4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X2B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X3B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X6B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P5M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P7M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1P4M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X2M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X3M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X4M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X2M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X3M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6B_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6M_A9TH (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X2M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X3M_A9TH (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P5M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P7M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1P4M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X2M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X3M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X4M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X6M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X8M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P5M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P7M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1P4M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X2M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X3M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X4M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X6M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X8M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nand (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P5M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P7M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1P4M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X2M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X3M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X4M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X6M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X8M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P5M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P7M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1P4M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X2M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X3M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X4M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X6M_A9TH (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P5M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P7M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1P4M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X2M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X3M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X4M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X6M_A9TH (Y,VDD, VSS, A, B, CN);
inout VDD, VSS;
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (out_temp, A, B, Cx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P5M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P7M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1P4M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X2M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X3M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X4M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X6M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P5M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P7M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1P4M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X2M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X3M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X4M_A9TH (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P5M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P7M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1P4M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X2M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X3M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X4M_A9TH (Y,VDD, VSS, A, B, C, DN);
inout VDD, VSS;
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (out_temp, A, B, C, Dx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4A_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P5M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P7M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1P4M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X2M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X3M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X4M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X6M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X8M_A9TH (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P5M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P7M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1P4M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X2M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X3M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X4M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X6M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X8M_A9TH (Y,VDD, VSS, A, BN);
inout VDD, VSS;
output Y;
input A, BN;

  not (Bx, BN);
  nor (out_temp, A, Bx);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8A_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P5M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P7M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1P4M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X2M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X3M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X4M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X6M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X8M_A9TH (Y,VDD, VSS, AN, BN, C);
inout VDD, VSS;
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4A_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P5M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P7M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1P4M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X2M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X3M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X4M_A9TH (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P5M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P7M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1P4M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X2M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X3M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X4M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X6M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X8M_A9TH (Y,VDD, VSS, A0N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (out_temp, A0N, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(out_temp, outB, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X8M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(out_temp, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X2M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X3M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X6M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X8M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X8M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X8M_A9TH (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X2M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X3M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X4M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X6M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X8M_A9TH (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X2M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X3M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X4M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X6M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X8M_A9TH (Y,VDD, VSS, A0, A1, B0N, B1N);
inout VDD, VSS;
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P5M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P7M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1P4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X2M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X3M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X4M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X6M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X8M_A9TH (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P5M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P7M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1P4M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X2M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X3M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X4M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X6M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X8M_A9TH (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P5M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P7M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1P4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X2M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X3M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X4M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X6M_A9TH (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8B_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X6M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X8M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X2M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X3M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X4M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X6M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X8M_A9TH (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P5M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P7M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1P4M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X2M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X3M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X4M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X6M_A9TH (Y,VDD, VSS, A, B, C, D, E, F);
inout VDD, VSS;
output Y;
input A, B, C, D, E, F;

  or (out_temp, A, B, C, D, E, F);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P5B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P6B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P7B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P8B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X11B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X13B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X16B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P2B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P4B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P7B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2P5B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3P5B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X4B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X5B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X6B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X7P5B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X9B_A9TH (ECK,VDD, VSS, CK, E, SEN);
inout VDD, VSS;
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat_PWR  I1 (n0, ovrd, CK, E, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P5B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P6B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P7B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P8B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X11B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X13B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X16B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P2B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P4B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P7B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2P5B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3P5B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X4B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X5B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X6B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X7P5B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X9B_A9TH (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1M_A9TH (RBL,VDD, VSS, RWL, WBL, WWL);
inout VDD, VSS;
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf_PWR  I0 (n0, WBL, WWL, wwn,  VDD, VSS, NOTIFIER);
   bufif1     I1 (rdbl_temp, n0, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1P4M_A9TH (RBL,VDD, VSS, RWL, WBL, WWL);
inout VDD, VSS;
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf_PWR  I0 (n0, WBL, WWL, wwn,  VDD, VSS, NOTIFIER);
   bufif1     I1 (rdbl_temp, n0, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X2M_A9TH (RBL,VDD, VSS, RWL, WBL, WWL);
inout VDD, VSS;
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf_PWR  I0 (n0, WBL, WWL, wwn,  VDD, VSS, NOTIFIER);
   bufif1     I1 (rdbl_temp, n0, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1M_A9TH (RBL,VDD, VSS, RWL, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(rdbl_temp, n1, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1P4M_A9TH (RBL,VDD, VSS, RWL, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(rdbl_temp, n1, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X2M_A9TH (RBL,VDD, VSS, RWL, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(rdbl_temp, n1, RWL);
  assign RBL = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL, WWL);
inout VDD, VSS;
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf_PWR  I3 (n0, WBL, WWL, WWLN,  VDD, VSS, NOTIFIER);
   bufif1     I4 (rdbl1_temp, n0, n2);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1     I5 (rdbl2_temp, n0, n3);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1P4M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL, WWL);
inout VDD, VSS;
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf_PWR  I3 (n0, WBL, WWL, WWLN,  VDD, VSS, NOTIFIER);
   bufif1     I4 (rdbl1_temp, n0, n2);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1     I5 (rdbl2_temp, n0, n3);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X2M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL, WWL);
inout VDD, VSS;
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf_PWR  I3 (n0, WBL, WWL, WWLN,  VDD, VSS, NOTIFIER);
   bufif1     I4 (rdbl1_temp, n0, n2);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1     I5 (rdbl2_temp, n0, n3);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (rdbl1_temp, n1, RWL1);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1 I6 (rdbl2_temp, n1, RWL2);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1P4M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (rdbl1_temp, n1, RWL1);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1 I6 (rdbl2_temp, n1, RWL2);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X2M_A9TH (RBL1, RBL2,VDD, VSS, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
inout VDD, VSS;
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2_PWR  I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, VDD, VSS, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (rdbl1_temp, n1, RWL1);
  assign RBL1 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   bufif1 I6 (rdbl2_temp, n1, RWL2);
  assign RBL2 = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFNQ_X1M_A9TH (Q,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X2M_A9TH (Q,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X3M_A9TH (Q,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X1M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X2M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X3M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X1M_A9TH (Q,VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X2M_A9TH (Q,VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X3M_A9TH (Q,VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X1M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X2M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X3M_A9TH (Q,VDD, VSS, CKN, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X1M_A9TH (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X2M_A9TH (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X3M_A9TH (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X1M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X2M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X3M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X4M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X1M_A9TH (QN,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X2M_A9TH (QN,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X3M_A9TH (QN,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X1M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X2M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X3M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X4M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X0P5M_A9TH (QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X1M_A9TH (QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X2M_A9TH (QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X3M_A9TH (QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X1M_A9TH (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X2M_A9TH (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X3M_A9TH (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X4M_A9TH (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X0P5M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X1M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X2M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X3M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X4M_A9TH (Q,VDD, VSS, CK, D, R, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X1M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X2M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X3M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X4M_A9TH (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module TIEHI_X1M_A9TH (Y,VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIEHI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO_X1M_A9TH (Y,VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIELO_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P5M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P7M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1P4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X2M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X3M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X4M_A9TH (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P5M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P7M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1P4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X2M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X3M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X4M_A9TH (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X4M_A9TH
`endcelldefine
`else

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X0P5M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X1M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X2M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQN_X3M_A9TH (QN, A, B, CK, SE, SI);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X0P5M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X1M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X2M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X3M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module A2SDFFQ_X4M_A9TH (Q, A, B, CK, SE, SI);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);

wire ENABLE_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_NOT_B_AND_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_NOT_SE_AND_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_NOT_SI ;
wire ENABLE_A_AND_B_AND_SE_AND_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SI ;
wire ENABLE_NOT_A_AND_B_AND_SI ;
wire ENABLE_A_AND_NOT_B_AND_SI ;
wire ENABLE_A_AND_B_AND_NOT_SI ;
wire ENABLE_NOT_A_AND_NOT_B_AND_SE ;
wire ENABLE_NOT_A_AND_B_AND_SE ;
wire ENABLE_A_AND_NOT_B_AND_SE ;
wire ENABLE_A_AND_B_AND_SE ;
assign ENABLE_B_AND_NOT_SE_AND_NOT_SI = (B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_B_AND_NOT_SE_AND_SI = (B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_NOT_SI = (A&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_SE_AND_SI = (A&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (!A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI = (!A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI = (!A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI = (!A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI = (!A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI = (!A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI = (!A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE_AND_SI = (!A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI = (A&!B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI = (A&!B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI = (A&!B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE_AND_SI = (A&!B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI = (A&B&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SE_AND_SI = (A&B&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_NOT_SI = (A&B&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE_AND_SI = (A&B&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SI = (!A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SI = (!A&B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SI = (A&!B&SI) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_NOT_SI = (A&B&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_NOT_B_AND_SE = (!A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_A_AND_B_AND_SE = (!A&B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_NOT_B_AND_SE = (A&!B&SE) ? 1'b1:1'b0;
assign ENABLE_A_AND_B_AND_SE = (A&B&SE) ? 1'b1:1'b0;

specify
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), posedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_B_AND_NOT_SE_AND_SI == 1'b1), negedge A, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), posedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_SE_AND_SI == 1'b1), negedge B, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_A_AND_B_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_NOT_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_A_AND_B_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (A==1'b0 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b0 && SI==1'b1 || A==1'b0 && B==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // A2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X1P4M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFCIN_X2M_A9TH ( CO, SUM, A, B, CIN);
output SUM, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (SUM, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X1P4M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X2M_A9TH ( CO, SUM, A, B, CI);
output SUM, CO;
input A, B, CI;
  xor I0(SUM, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1P4M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X2M_A9TH ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1P4M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X2M_A9TH ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X11M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X11M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X8M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X6M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X8M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X8M_A9TH
`endcelldefine
module ANTENNA1_A9TH (A);
input A;


specify

endspecify
endmodule // ANTENNA1_A9TH
`timescale 1ns/1ps
`celldefine
module AO1B2_X0P5M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X0P7M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X1P4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X2M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X3M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO1B2_X6M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P5M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X0P7M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1P4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X2M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X3M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P5M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P7M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1P4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X2M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X3M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P5M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P7M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X1P4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X2M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X3M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X6M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X8M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P5M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P7M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X1P4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X2M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X3M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X6M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X8M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P5M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P7M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1P4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X2M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X3M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X6M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P5M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X0P7M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1P4M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X2M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X3M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X4M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X6M_A9TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X11M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X16M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X2M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X3M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X4M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X6M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENC_X8M_A9TH (AN, SN, X2, M0, M1, M2);
output SN, AN, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (SN, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (AN, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => AN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => SN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENC_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X0P7M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN, nPP);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN, nPP);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X1P4M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN, nPP);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXIT_X2M_A9TH (PPN, AN, D0, D1, SN, X2);
output PPN;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (nPP, X2, AN, SN, D1, D0);
  not  I1 (PPN, nPP);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PPN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PPN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXIT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X0P7M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (PP, X2, AN, SN, D1, D0);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (PP, X2, AN, SN, D1, D0);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X1P4M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (PP, X2, AN, SN, D1, D0);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXT_X2M_A9TH (PP, AN, D0, D1, SN, X2);
output PP;
input X2, AN, SN, D1, D0;

  udp_bmx I0 (PP, X2, AN, SN, D1, D0);



specify
if (D0==1'b0 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b0 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b0)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && SN==1'b1 && X2==1'b1)
(AN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(posedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1)
(negedge D0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(posedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1)
(negedge D1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b0 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && X2==1'b1)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && X2==1'b0)
(SN => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b0 && D1==1'b1 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b1 && D1==1'b0 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b0 && D0==1'b1 && D1==1'b0 && SN==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (AN==1'b1 && D0==1'b0 && D1==1'b1 && SN==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXT_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P7M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X0P8M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X11M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X13M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X16M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P2M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P4M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X1P7M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X2P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X3P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X4M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X6M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X7P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFH_X9M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFH_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X11M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X16M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X1P4M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X2M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X3M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X4M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X6M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFZ_X8M_A9TH ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFZ_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P7M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X0P8M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X11M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X13M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P2M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P4M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X1P7M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X7P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X9M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X1P4M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCIN_X2M_A9TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCIN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X1P4M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENCON_X2M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENCON_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1P4M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X2M_A9TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1P4M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X2M_A9TH ( CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (CO, t5, t6, t7);



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X1P4M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (CO, t5, t6, t7);



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42_X2M_A9TH (CO, ICO, SUM, A, B, C, D, ICI);
output SUM, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor  I7 (SUM, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (CO, t5, t6, t7);



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => SUM) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFNQ_X1M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X2M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNQ_X3M_A9TH (Q, CKN, D);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X1M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X2M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRPQ_X3M_A9TH (Q, CKN, D, R, SN);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_NOT_D ;
wire ENABLE_NOT_CKN_AND_D ;
wire ENABLE_CKN_AND_NOT_D ;
wire ENABLE_CKN_AND_D ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CKN_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SN = (!CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SN = (!CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SN = (CKN&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SN = (CKN&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D = (!CKN&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D = (!CKN&D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D = (CKN&!D) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D = (CKN&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R = (!CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R = (!CKN&D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R = (CKN&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R = (CKN&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X0P5M_A9TH (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X1M_A9TH (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X2M_A9TH (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X3M_A9TH (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X0P5M_A9TH (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X1M_A9TH (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X2M_A9TH (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X3M_A9TH (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X4M_A9TH (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X0P5M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X1M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X2M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQN_X3M_A9TH (QN, CK, D, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFRPQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X0P5M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X1M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X2M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X3M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRPQ_X4M_A9TH (Q, CK, D, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X0P5M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X1M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X2M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQN_X3M_A9TH (QN, CK, D, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  not     I2 (QN, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSQN_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X0P5M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X1M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X2M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X3M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X4M_A9TH (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X0P5M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X0P5M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X1M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X1M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X2M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X2M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X3M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X3M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRPQ_X4M_A9TH (Q, CK, D, R, SN);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SN ;
wire ENABLE_NOT_R_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SN ;
wire ENABLE_CK_AND_D_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_NOT_D ;
wire ENABLE_NOT_CK_AND_D ;
wire ENABLE_CK_AND_NOT_D ;
wire ENABLE_CK_AND_D ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R ;
wire ENABLE_CK_AND_D_AND_NOT_R ;
assign ENABLE_NOT_D_AND_NOT_R_AND_SN = (!D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SN = (D&!R&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_SN = (!R&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SN = (!CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SN = (!CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SN = (CK&!D&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SN = (CK&D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D = (!CK&!D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D = (!CK&D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D = (CK&!D) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D = (CK&D) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R = (!CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R = (!CK&D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R = (CK&!D&!R) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R = (CK&D&!R) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRPQ_X4M_A9TH
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY2_X0P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X1M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X0P5M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X1M_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S2_X1B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S4_X1B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S4_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S6_X1B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S6_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLYCLK8S8_X1B_A9TH ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLYCLK8S8_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ENDCAPTIE3_A9TH;

endmodule //ENDCAPTIE3_A9TH

`endcelldefine
`timescale 1ns/1ps
`celldefine
module ESDFFQN_X0P5M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X1M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X2M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQN_X3M_A9TH (QN, CK, D, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQN_X3M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X0P5M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X0P5M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X1M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X1M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X2M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X2M_A9TH
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ESDFFQ_X3M_A9TH (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_E_AND_SE_AND_SI ;
wire ENABLE_E_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_E_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SI ;
wire ENABLE_NOT_D_AND_E_AND_SI ;
wire ENABLE_D_AND_NOT_E_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_E_AND_SI ;
wire ENABLE_D_AND_E_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_E_AND_SE ;
wire ENABLE_NOT_D_AND_E_AND_SE ;
wire ENABLE_D_AND_NOT_E_AND_SE ;
wire ENABLE_D_AND_E_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI = (!D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI = (!D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI = (!D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI = (!D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI = (!D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE_AND_SI = (!D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI = (D&!E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE_AND_SI = (D&!E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI = (D&E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SE_AND_SI = (D&E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_NOT_SI = (D&E&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE_AND_SI = (D&E&SE&SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_NOT_SI = (E&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE_AND_SI = (E&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI = (!D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SI = (!D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SI = (!D&E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_NOT_SI = (D&!E&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SI = (D&!E&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_NOT_SI = (D&E&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_E_AND_SE = (!D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_E_AND_SE = (!D&E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_E_AND_SE = (D&!E&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_E_AND_SE = (D&E&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_E_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ESDFFQ_X3M_A9TH
`endcelldefine


module FILL128_A9TH;

endmodule //FILL128_A9TH


module FILL16_A9TH;

endmodule //FILL16_A9TH


module FILL1_A9TH;

endmodule //FILL1_A9TH


module FILL2_A9TH;

endmodule //FILL2_A9TH


module FILL32_A9TH;

endmodule //FILL32_A9TH


module FILL4_A9TH;

endmodule //FILL4_A9TH


module FILL64_A9TH;

endmodule //FILL64_A9TH


module FILL8_A9TH;

endmodule //FILL8_A9TH


module FILLCAP128_A9TH;


specify

endspecify
endmodule // FILLCAP128_A9TH

module FILLCAP16_A9TH;


specify

endspecify
endmodule // FILLCAP16_A9TH

module FILLCAP32_A9TH;


specify

endspecify
endmodule // FILLCAP32_A9TH

module FILLCAP4_A9TH;


specify

endspecify
endmodule // FILLCAP4_A9TH

module FILLCAP64_A9TH;


specify

endspecify
endmodule // FILLCAP64_A9TH

module FILLCAP8_A9TH;


specify

endspecify
endmodule // FILLCAP8_A9TH

module FILLSGCAP128_A9TH;


specify

endspecify
endmodule // FILLSGCAP128_A9TH

module FILLSGCAP16_A9TH;


specify

endspecify
endmodule // FILLSGCAP16_A9TH

module FILLSGCAP32_A9TH;


specify

endspecify
endmodule // FILLSGCAP32_A9TH

module FILLSGCAP4_A9TH;


specify

endspecify
endmodule // FILLSGCAP4_A9TH

module FILLSGCAP64_A9TH;


specify

endspecify
endmodule // FILLSGCAP64_A9TH

module FILLSGCAP8_A9TH;


specify

endspecify
endmodule // FILLSGCAP8_A9TH

module FILLTIE128_A9TH;

endmodule //FILLTIE128_A9TH


module FILLTIE16_A9TH;

endmodule //FILLTIE16_A9TH


module FILLTIE32_A9TH;

endmodule //FILLTIE32_A9TH


module FILLTIE3_A9TH;

endmodule //FILLTIE3_A9TH


module FILLTIE4_A9TH;

endmodule //FILLTIE4_A9TH


module FILLTIE64_A9TH;

endmodule //FILLTIE64_A9TH


module FILLTIE8_A9TH;

endmodule //FILLTIE8_A9TH


`timescale 1ns/1ps
`celldefine
module FRICG_X0P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P6B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P7B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X0P8B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X11B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X13B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X16B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P2B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P4B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X1P7B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X2P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X3P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X4B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X6B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X7P5B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FRICG_X9B_A9TH ( ECK, CK );
output ECK;
input CK;

  buf I0(ECK, CK);



specify
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // FRICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P6M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P7M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P8M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X11M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X13M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X13M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P2M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P4M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1P7M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2P5M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3P5M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X7P5M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X7P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9B_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X9M_A9TH ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X9M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X0P5M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X1M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X2M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X3M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQN_X4M_A9TH (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X0P5M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X1M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X2M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNQ_X3M_A9TH (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATNQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X0P5M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X1M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X2M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X3M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRPQN_X4M_A9TH (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X0P5M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X1M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X2M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNRQ_X3M_A9TH (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X0P5M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X1M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X2M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSPQ_X3M_A9TH (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATNSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X0P5M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X1M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X2M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X3M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATNSQN_X4M_A9TH (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_GN ;
wire ENABLE_D_AND_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_GN = (!D&GN) ? 1'b1:1'b0;
assign ENABLE_D_AND_GN = (D&GN) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_GN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATNSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X0P5M_A9TH (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X1M_A9TH (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X2M_A9TH (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X3M_A9TH (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQN_X4M_A9TH (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X0P5M_A9TH (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X1M_A9TH (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X2M_A9TH (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATQ_X3M_A9TH (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // LATQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X0P5M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X1M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X2M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X3M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRPQN_X4M_A9TH (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_NOT_R ;
wire ENABLE_NOT_D_AND_NOT_R ;
wire ENABLE_D_AND_NOT_R ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R = (!D&!R) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R = (D&!R) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_R == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_R == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge R, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(R => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRPQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X0P5M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X1M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X2M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATRQ_X3M_A9TH (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_D_AND_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN = (D&RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge RN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // LATRQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X0P5M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X1M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X2M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSPQ_X3M_A9TH (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not  I3(clk,G);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_D_AND_NOT_S ;
wire ENABLE_D_AND_NOT_S ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_S = (!D&!S) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_S = (D&!S) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_NOT_S == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_NOT_S == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(negedge S, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge S &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1)
(S => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // LATSPQ_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X0P5M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X1M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X2M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X3M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module LATSQN_X4M_A9TH (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_D_AND_NOT_G ;
wire ENABLE_D_AND_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SN = (!D&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_G = (!D&!G) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_G = (D&!G) ? 1'b1:1'b0;

specify
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_NOT_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_D_AND_NOT_G == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // LATSQN_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X0P5M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X1M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X2M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQN_X3M_A9TH (QN, CK, D0, D1, S0, SE, SI);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X0P5M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X1M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X2M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X3M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module M2SDFFQ_X4M_A9TH (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI ;
wire ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE ;
wire ENABLE_D0_AND_D1_AND_S0_AND_SE ;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (!D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (!D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (!D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (!D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (!D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI = (!D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&!D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&!D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&!D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&!D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&!D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI = (D0&!D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D0&D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI = (D0&D1&!S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI = (D0&D1&!S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&D1&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI = (D0&D1&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI = (D0&D1&S0&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI = (D0&D1&S0&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (!D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (!D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI = (D1&!S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI = (D1&!S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (!D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI = (!D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI = (D0&S0&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI = (D0&S0&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI = (!D0&D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI = (!D0&D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI = (D0&!D1&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI = (D0&!D1&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI = (!D0&!D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI = (!D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI = (!D0&D1&!S0&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI = (!D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI = (D0&!D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI = (D0&!D1&S0&SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI = (D0&D1&!S0&!SI) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI = (D0&D1&S0&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (!D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE = (!D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE = (!D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE = (!D0&D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE = (D0&!D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE = (D0&!D1&S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE = (D0&D1&!S0&SE) ? 1'b1:1'b0;
assign ENABLE_D0_AND_D1_AND_S0_AND_SE = (D0&D1&S0&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_S0_AND_NOT_SE_AND_SI == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_SE_AND_SI == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_NOT_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_NOT_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D0_AND_D1_AND_S0_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // M2SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module MX2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X8B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXGL2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXGL2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P5M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X0P7M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X1P4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X2M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X3M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT2_X4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P5M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X0P7M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X1P4M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X2M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXIT4_X3M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXIT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P5M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X0P7M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X1P4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X2M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X3M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X4M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6B_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT2_X6M_A9TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P5M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X0P7M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X1P4M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X2M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXT4_X3M_A9TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXT4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P5M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X0P7M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1P4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X2M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X3M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X6M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X8M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P5M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P7M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X1P4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X2M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X3M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X6M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X8M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8A_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P5M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P7M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X1P4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X2M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X3M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X6M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X8M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P5M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X0P7M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1P4M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X2M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X3M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X4M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X6M_A9TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P5M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X0P7M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X1P4M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X2M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X3M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X4M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XXB_X6M_A9TH (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XXB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P5M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X0P7M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1P4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X2M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X3M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X6M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P5M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X0P7M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1P4M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X2M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X3M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X4M_A9TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P5M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X0P7M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X1P4M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X2M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X3M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XXXB_X4M_A9TH (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(DN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XXXB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4A_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P5M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X0P7M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1P4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X2M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X3M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X4M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X6M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X8M_A9TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P5M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P7M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X1P4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X2M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X3M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X4M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X6M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X8M_A9TH (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8A_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P5M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P7M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X1P4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X2M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X3M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X4M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X6M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X8M_A9TH (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P5A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P7A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1P4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X3A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4A_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4A_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P5M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X0P7M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1P4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X2M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X3M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X4M_A9TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P5M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P7M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X1P4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X2M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X3M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X4M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X6M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X8M_A9TH (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X6M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not I0(outB, B0N);
  or  I1(outA, A0, A1);
  and I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P5M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P7M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1P4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X2M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X3M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X4M_A9TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P5M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P7M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1P4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X2M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X3M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X4M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X6M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X8M_A9TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P5M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P7M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1P4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X2M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X3M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X4M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X6M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X8M_A9TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P5M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X0P7M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1P4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X2M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X3M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X4M_A9TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P5M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P7M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1P4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X2M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X3M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X4M_A9TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P5M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P7M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X1P4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X2M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X3M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X4M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X6M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X8M_A9TH (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P5M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P7M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1P4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X2M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X3M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X4M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X6M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X8M_A9TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P5M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X0P7M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X1P4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X2M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X3M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X4M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X6M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2XB1_X8M_A9TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2XB1_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P5M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P7M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1P4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X2M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X3M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X4M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X6M_A9TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X11M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X11M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8B_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8M_A9TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X6M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X8M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P5M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X0P7M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1P4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X2M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X3M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X4M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X6M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X8M_A9TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X8M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P5M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X0P7M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X1P4M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X2M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X3M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X4M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR6_X6M_A9TH (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(E => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(F => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR6_X6M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P6B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P7B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X0P8B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X11B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X13B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X16B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P2B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P4B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X1P7B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X2P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X3P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X4B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X6B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X7P5B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module POSTICG_X9B_A9TH (ECK, CK, E, SEN);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_SEN ;
wire ENABLE_E_AND_SEN ;
wire ENABLE_SEN ;
wire ENABLE_NOT_E ;
wire ENABLE_CK_AND_NOT_E ;
wire ENABLE_CK_AND_E ;
assign ENABLE_NOT_E_AND_SEN = (!E&SEN) ? 1'b1:1'b0;
assign ENABLE_E_AND_SEN = (E&SEN) ? 1'b1:1'b0;
assign ENABLE_SEN = (SEN) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_E = (CK&!E) ? 1'b1:1'b0;
assign ENABLE_CK_AND_E = (CK&E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SEN==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SEN==1'b1)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SEN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SEN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SEN, posedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SEN &&& (ENABLE_CK_AND_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (E==1'b0)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (E==1'b1)
(negedge SEN *> (ECK +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // POSTICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P6B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P7B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X0P8B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X0P8B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X11B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X11B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X13B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X13B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X16B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X16B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P2B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P4B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X1P7B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X1P7B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X2B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X2P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X2P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X3B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X3P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X3P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X4B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X4B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X6B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X6B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X7P5B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X7P5B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module PREICG_X9B_A9TH (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_NOT_E_AND_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_E_AND_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E_AND_SE = (!E&SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_SE = (E&SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_AND_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // PREICG_X9B_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X1P4M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WS_X2M_A9TH (RBL, RWL, WBL, WWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn,  NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);





wire ENABLE_RWL ;
wire ENABLE_RWL_AND_NOT_WBL ;
wire ENABLE_RWL_AND_WBL ;
assign ENABLE_RWL = (RWL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL = (RWL&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL = (RWL&WBL) ? 1'b1:1'b0;

specify
(WBL => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b0 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL==1'b1 && WWL==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WWL==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge WWL => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(RBL, n1, RWL);





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X1P4M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(RBL, n1, RWL);





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R2WS_X2M_A9TH (RBL, RWL, WBL1, WBL2, WWL1, WWL2);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1   I5(RBL, n1, RWL);





wire ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 = (RWL&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (WBL2==1'b0)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(WBL1 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(WBL2 => RBL) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL => RBL ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL => RBL ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (WBL2==1'b0)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL2==1'b1)
(posedge WWL1 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b0)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WBL1==1'b1)
(posedge WWL2 => (RBL:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X1P4M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WS_X2M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL, WWL);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN,  NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2 ;
wire ENABLE_RWL1_AND_RWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL ;
assign ENABLE_NOT_RWL1_AND_RWL2 = (!RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2 = (RWL1&!RWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2 = (RWL1&RWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL = (!RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL = (!RWL1&RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL = (RWL1&!RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL = (RWL1&!RWL2&WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL = (RWL1&RWL2&!WBL) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL = (RWL1&RWL2&WBL) ? 1'b1:1'b0;

specify
if (RWL2==1'b0)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(WBL => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(WBL => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WWL==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b0 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL==1'b1 && WWL==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WWL==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), posedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL &&& (ENABLE_RWL1_AND_RWL2 == 1'b1), negedge WBL, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL &&& (ENABLE_RWL1_AND_RWL2_AND_WBL == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1)
(posedge WWL => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1)
(posedge WWL => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (RBL1, n1, RWL1);
   bufif1 I6 (RBL2, n1, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X1P4M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (RBL1, n1, RWL1);
   bufif1 I6 (RBL2, n1, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R2WS_X2M_A9TH (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   not I1 (WBL1_not, WBL1);
   not I2 (WBL2_not, WBL2);
   udp_tlatrf2 I3 (n0, WBL1_not, WWL1, WBL2_not, WWL2, NOTIFIER);
   not I4 (n1, n0);
   bufif1 I5 (RBL1, n1, RWL1);
   bufif1 I6 (RBL2, n1, RWL2);





wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 ;
wire ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 ;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (!RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&!RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&!WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&!WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 = (RWL1&RWL2&WBL1&WBL2&!WWL2) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (!RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&!RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&!WBL1&WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&!WBL2&!WWL1) ? 1'b1:1'b0;
assign ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 = (RWL1&RWL2&WBL1&WBL2&!WWL1) ? 1'b1:1'b0;

specify
if (RWL2==1'b0 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(WBL1 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(WBL2 => RBL1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(WBL1 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(WBL2 => RBL2) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL2==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL1 => RBL1 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL2==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL1 => RBL1 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b0 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b0 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b0 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY,0);
if (RWL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b0)
( RWL2 => RBL2 ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b0 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WWL1==1'b0 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1 && WBL2==1'b1 && WWL1==1'b1 && WWL2==1'b1 || RWL1==1'b1 && WBL1==1'b0 && WBL2==1'b0 && WWL1==1'b1 && WWL2==1'b1)
( RWL2 => RBL2 ) = (0, 0, 0,`ARM_PROP_DELAY, 0,`ARM_PROP_DELAY);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), posedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL2_AND_NOT_WWL2 == 1'b1), negedge WBL1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), posedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WWL1 == 1'b1), negedge WBL2, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL1 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL2 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_NOT_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_NOT_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_NOT_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_NOT_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge WWL2 &&& (ENABLE_RWL1_AND_RWL2_AND_WBL1_AND_WBL2_AND_NOT_WWL1 == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (RWL2==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL2==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL1:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b0)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL2==1'b1)
(posedge WWL1 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b0 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b0)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RWL1==1'b1 && WBL1==1'b1)
(posedge WWL2 => (RBL2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R2WS_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFNQ_X1M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X2M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNQ_X3M_A9TH (Q, CKN, D, SE, SI);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X1M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X2M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRPQ_X3M_A9TH (Q, CKN, D, R, SE, SI);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X1M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X2M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSQ_X3M_A9TH (Q, CKN, D, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFNSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X1M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X2M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQ_X3M_A9TH (Q, CKN, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN = (!CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CKN&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CKN&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CKN&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CKN&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN = (CKN&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (!CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (!CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI = (!CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI = (!CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI = (!CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI = (!CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI = (CKN&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI = (CKN&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI = (CKN&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI = (CKN&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI = (CKN&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI = (CKN&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_SE_AND_SI = (CKN&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CKN&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CKN&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CKN&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CKN&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CKN&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI = (CKN&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, negedge CKN &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CKN_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CKN_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X0P5M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X1M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X2M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X3M_A9TH (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X0P5M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X1M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X2M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X3M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X4M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X0P5M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X1M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X2M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQN_X3M_A9TH (QN, CK, D, R, SE, SI);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFRPQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X0P5M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X1M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X2M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X3M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRPQ_X4M_A9TH (Q, CK, D, R, SE, SI);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE ;
wire ENABLE_D_AND_NOT_R_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI = (D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI = (D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI = (!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI = (!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI = (!D&!R&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI = (D&!R&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE = (!D&!R&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE = (D&!R&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X0P5M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X1M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X2M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQN_X3M_A9TH (QN, CK, D, SE, SI, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSQN_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X0P5M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X1M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X2M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X3M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X4M_A9TH (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SN ;
wire ENABLE_D_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI_AND_SN = (D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI_AND_SN = (!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI_AND_SN = (!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI_AND_SN = (!D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN = (D&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SN = (!D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SN = (D&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X0P5M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X0P5M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X1M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X2M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X3M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRPQ_X4M_A9TH (Q, CK, D, R, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI ;
wire ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI ;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (!D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (!D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (D&!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN = (D&!R&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN = (D&!R&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN = (!R&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN = (!R&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI_AND_SN = (!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI_AND_SN = (D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI_AND_SN = (D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (!CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (!CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (!CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (!CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN = (!CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&!D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN = (CK&!D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN = (CK&!D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN = (CK&!D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN = (CK&D&!SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN = (CK&D&!SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN = (CK&D&SE&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN = (CK&D&SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN = (!D&!R&SI&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN = (D&!R&!SI&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN = (!D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_SN = (D&!R&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI = (D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (!CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (!CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI = (!CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (!CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI = (!CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI = (!CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_SE_AND_SI = (!CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI = (CK&!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI = (CK&!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI = (CK&!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_SE_AND_SI = (CK&!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI = (CK&D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_SE_AND_SI = (CK&D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_NOT_SI = (CK&D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_SE_AND_SI = (CK&D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (!CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (!CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (!CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (!CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (!CK&D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&!D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&!D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&!D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI = (CK&!D&!R&SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI = (CK&D&!R&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI = (CK&D&!R&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI = (CK&D&!R&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI = (CK&D&!R&SE&SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_R_AND_NOT_SE_AND_SI_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(negedge R, posedge CK &&& (ENABLE_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_NOT_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_NOT_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_NOT_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_NOT_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_NOT_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R &&& (ENABLE_CK_AND_D_AND_SE_AND_SI == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_NOT_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge SN &&& (ENABLE_CK_AND_D_AND_NOT_R_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(posedge R *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && R==1'b1 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRPQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X1M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X1M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X2M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X2M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X3M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X3M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFYQ_X4M_A9TH (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SE_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE_AND_SI ;
wire ENABLE_D_AND_NOT_SE_AND_NOT_SI ;
wire ENABLE_D_AND_NOT_SE_AND_SI ;
wire ENABLE_D_AND_SE_AND_NOT_SI ;
wire ENABLE_D_AND_SE_AND_SI ;
wire ENABLE_NOT_SE_AND_NOT_SI ;
wire ENABLE_NOT_SE_AND_SI ;
wire ENABLE_NOT_D_AND_SI ;
wire ENABLE_D_AND_NOT_SI ;
wire ENABLE_NOT_D_AND_SE ;
wire ENABLE_D_AND_SE ;
assign ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI = (!D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_AND_SI = (!D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_NOT_SI = (!D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE_AND_SI = (!D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_NOT_SI = (D&!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SI = (D&!SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_NOT_SI = (D&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE_AND_SI = (D&SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_NOT_SI = (!SE&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SI = (!SE&SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SI = (!D&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI = (D&!SI) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_SE = (!D&SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_SE = (D&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_NOT_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(posedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_D_AND_SE_AND_SI == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_NOT_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SI == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFYQ_X4M_A9TH
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module TIEHI_X1M_A9TH (Y);
output Y;

  buf I0(Y, 1'b1);


specify

endspecify
endmodule // TIEHI_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO_X1M_A9TH (Y);
output Y;

  buf I0(Y, 1'b0);


specify

endspecify
endmodule // TIELO_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P5M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P7M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1P4M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X2M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X3M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X4M_A9TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P5M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X0P5M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P7M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X0P7M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1P4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1P4M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X2M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X2M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X3M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X3M_A9TH
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X4M_A9TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X4M_A9TH
`endcelldefine
`endif
`endif
